library verilog;
use verilog.vl_types.all;
entity rw_manager_core is
    generic(
        AVL_DATA_WIDTH  : string  := "";
        AVL_ADDRESS_WIDTH: string  := "";
        MEM_DQ_WIDTH    : string  := "";
        MEM_DM_WIDTH    : string  := "";
        MEM_ODT_WIDTH   : string  := "";
        MEM_NUMBER_OF_RANKS: string  := "";
        AC_ODT_BIT      : string  := "";
        AC_BUS_WIDTH    : string  := "";
        AC_MASKED_BUS_WIDTH: string  := "";
        MASK_WIDTH      : string  := "";
        AFI_RATIO       : string  := "";
        MEM_READ_DQS_WIDTH: string  := "";
        MEM_WRITE_DQS_WIDTH: string  := "";
        DEBUG_READ_DI_WIDTH: string  := "";
        DEBUG_WRITE_TO_READ_RATIO_2_EXPONENT: string  := "";
        DEBUG_WRITE_TO_READ_RATIO: string  := "";
        MAX_DI_BUFFER_WORDS_LOG_2: string  := "";
        RATE            : string  := "";
        HCX_COMPAT_MODE : integer := 0;
        DEVICE_FAMILY   : string  := "";
        AC_ROM_INIT_FILE_NAME: string  := "AC_ROM.hex";
        INST_ROM_INIT_FILE_NAME: string  := "inst_ROM.hex";
        USE_ALL_AFI_PHASES_FOR_COMMAND_ISSUE: integer := 0
    );
    port(
        avl_clk         : in     vl_logic;
        avl_reset_n     : in     vl_logic;
        avl_address     : in     vl_logic_vector;
        avl_readdata    : out    vl_logic_vector;
        avl_writedata   : in     vl_logic_vector;
        afi_clk         : in     vl_logic;
        afi_reset_n     : in     vl_logic;
        afi_wdata       : out    vl_logic_vector;
        afi_dm          : out    vl_logic_vector;
        afi_rdata       : in     vl_logic_vector;
        afi_rdata_valid : in     vl_logic;
        afi_rrank       : out    vl_logic_vector;
        afi_wrank       : out    vl_logic_vector;
        afi_odt         : out    vl_logic_vector;
        ac_masked_bus   : out    vl_logic_vector;
        ac_bus          : out    vl_logic_vector;
        cmd_read        : in     vl_logic;
        cmd_write       : in     vl_logic;
        cmd_done        : out    vl_logic;
        csr_clk         : in     vl_logic;
        csr_ena         : in     vl_logic;
        csr_dout_phy    : in     vl_logic;
        csr_dout        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AVL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AVL_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_NUMBER_OF_RANKS : constant is 1;
    attribute mti_svvh_generic_type of AC_ODT_BIT : constant is 1;
    attribute mti_svvh_generic_type of AC_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AC_MASKED_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MASK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATIO : constant is 1;
    attribute mti_svvh_generic_type of MEM_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_READ_DI_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_WRITE_TO_READ_RATIO_2_EXPONENT : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_WRITE_TO_READ_RATIO : constant is 1;
    attribute mti_svvh_generic_type of MAX_DI_BUFFER_WORDS_LOG_2 : constant is 1;
    attribute mti_svvh_generic_type of RATE : constant is 1;
    attribute mti_svvh_generic_type of HCX_COMPAT_MODE : constant is 1;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of AC_ROM_INIT_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of INST_ROM_INIT_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of USE_ALL_AFI_PHASES_FOR_COMMAND_ISSUE : constant is 1;
end rw_manager_core;
