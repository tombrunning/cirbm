library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_axi_st_converter is
    generic(
        AXI_ID_WIDTH    : integer := 4;
        AXI_ADDR_WIDTH  : integer := 32;
        AXI_LEN_WIDTH   : integer := 4;
        AXI_SIZE_WIDTH  : integer := 3;
        AXI_BURST_WIDTH : integer := 2;
        AXI_LOCK_WIDTH  : integer := 2;
        AXI_CACHE_WIDTH : integer := 4;
        AXI_PROT_WIDTH  : integer := 3;
        AXI_DATA_WIDTH  : integer := 32;
        AXI_RESP_WIDTH  : integer := 4;
        ST_ADDR_WIDTH   : integer := 32;
        ST_SIZE_WIDTH   : integer := 5;
        ST_ID_WIDTH     : integer := 4;
        ST_DATA_WIDTH   : integer := 32;
        COMMAND_ARB_TYPE: string  := "ROUND_ROBIN";
        REGISTERED      : integer := 1
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        awid            : in     vl_logic_vector;
        awaddr          : in     vl_logic_vector;
        awlen           : in     vl_logic_vector;
        awsize          : in     vl_logic_vector;
        awburst         : in     vl_logic_vector;
        awlock          : in     vl_logic_vector;
        awcache         : in     vl_logic_vector;
        awprot          : in     vl_logic_vector;
        awvalid         : in     vl_logic;
        awready         : out    vl_logic;
        wid             : in     vl_logic_vector;
        wdata           : in     vl_logic_vector;
        wstrb           : in     vl_logic_vector;
        wlast           : in     vl_logic;
        wvalid          : in     vl_logic;
        wready          : out    vl_logic;
        bid             : out    vl_logic_vector;
        bresp           : out    vl_logic_vector;
        bvalid          : out    vl_logic;
        bready          : in     vl_logic;
        arid            : in     vl_logic_vector;
        araddr          : in     vl_logic_vector;
        arlen           : in     vl_logic_vector;
        arsize          : in     vl_logic_vector;
        arburst         : in     vl_logic_vector;
        arlock          : in     vl_logic_vector;
        arcache         : in     vl_logic_vector;
        arprot          : in     vl_logic_vector;
        arvalid         : in     vl_logic;
        arready         : out    vl_logic;
        rid             : out    vl_logic_vector;
        rdata           : out    vl_logic_vector;
        rresp           : out    vl_logic_vector;
        rlast           : out    vl_logic;
        rvalid          : out    vl_logic;
        rready          : in     vl_logic;
        itf_cmd_ready   : in     vl_logic;
        itf_cmd_valid   : out    vl_logic;
        itf_cmd         : out    vl_logic;
        itf_cmd_address : out    vl_logic_vector;
        itf_cmd_burstlen: out    vl_logic_vector;
        itf_cmd_id      : out    vl_logic_vector;
        itf_cmd_priority: out    vl_logic;
        itf_cmd_autoprecharge: out    vl_logic;
        itf_cmd_multicast: out    vl_logic;
        itf_wr_data_ready: in     vl_logic;
        itf_wr_data_valid: out    vl_logic;
        itf_wr_data     : out    vl_logic_vector;
        itf_wr_data_byte_en: out    vl_logic_vector;
        itf_wr_data_begin: out    vl_logic;
        itf_wr_data_last: out    vl_logic;
        itf_wr_data_id  : out    vl_logic_vector;
        itf_rd_data_ready: out    vl_logic;
        itf_rd_data_valid: in     vl_logic;
        itf_rd_data     : in     vl_logic_vector;
        itf_rd_data_error: in     vl_logic;
        itf_rd_data_begin: in     vl_logic;
        itf_rd_data_last: in     vl_logic;
        itf_rd_data_id  : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AXI_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_LEN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_BURST_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_LOCK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_CACHE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_PROT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AXI_RESP_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ST_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ST_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ST_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ST_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of COMMAND_ARB_TYPE : constant is 1;
    attribute mti_svvh_generic_type of REGISTERED : constant is 1;
end alt_mem_ddrx_axi_st_converter;
