library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_csr is
    generic(
        DWIDTH_RATIO    : integer := 2;
        CTL_CSR_ENABLED : integer := 1;
        CTL_ECC_CSR_ENABLED: integer := 1;
        CTL_CSR_READ_ONLY: integer := 0;
        CTL_ECC_CSR_READ_ONLY: integer := 0;
        CFG_AVALON_ADDR_WIDTH: integer := 8;
        CFG_AVALON_DATA_WIDTH: integer := 32;
        MEM_IF_CLK_PAIR_COUNT: integer := 1;
        MEM_IF_DQS_WIDTH: integer := 72;
        \CFG_CS_ADDR_WIDTH\: integer := 1;
        \CFG_ROW_ADDR_WIDTH\: integer := 13;
        \CFG_COL_ADDR_WIDTH\: integer := 10;
        \CFG_BANK_ADDR_WIDTH\: integer := 3;
        \CFG_ENABLE_ECC\: integer := 1;
        \CFG_ENABLE_AUTO_CORR\: integer := 1;
        \CFG_REGDIMM_ENABLE\: integer := 0;
        CAS_WR_LAT_BUS_WIDTH: integer := 4;
        ADD_LAT_BUS_WIDTH: integer := 4;
        TCL_BUS_WIDTH   : integer := 4;
        BL_BUS_WIDTH    : integer := 5;
        TRRD_BUS_WIDTH  : integer := 4;
        TFAW_BUS_WIDTH  : integer := 6;
        TRFC_BUS_WIDTH  : integer := 8;
        TREFI_BUS_WIDTH : integer := 13;
        TRCD_BUS_WIDTH  : integer := 4;
        TRP_BUS_WIDTH   : integer := 4;
        TWR_BUS_WIDTH   : integer := 4;
        TWTR_BUS_WIDTH  : integer := 4;
        TRTP_BUS_WIDTH  : integer := 4;
        TRAS_BUS_WIDTH  : integer := 5;
        TRC_BUS_WIDTH   : integer := 6;
        AUTO_PD_BUS_WIDTH: integer := 16;
        STARVE_LIMIT_BUS_WIDTH: integer := 8;
        \CFG_CAS_WR_LAT\: integer := 0;
        \CFG_ADD_LAT\   : integer := 0;
        \CFG_TCL\       : integer := 0;
        \CFG_BURST_LENGTH\: integer := 0;
        \CFG_TRRD\      : integer := 0;
        \CFG_TFAW\      : integer := 0;
        \CFG_TRFC\      : integer := 0;
        \CFG_TREFI\     : integer := 0;
        \CFG_TRCD\      : integer := 0;
        \CFG_TRP\       : integer := 0;
        \CFG_TWR\       : integer := 0;
        \CFG_TWTR\      : integer := 0;
        \CFG_TRTP\      : integer := 0;
        \CFG_TRAS\      : integer := 0;
        \CFG_TRC\       : integer := 0;
        \CFG_AUTO_PD_CYCLES\: integer := 0;
        \CFG_ADDR_ORDER\: integer := 1;
        \CFG_REORDER_DATA\: integer := 0;
        \CFG_STARVE_LIMIT\: integer := 0;
        MEM_IF_CSR_COL_WIDTH: integer := 5;
        MEM_IF_CSR_ROW_WIDTH: integer := 5;
        MEM_IF_CSR_BANK_WIDTH: integer := 3;
        MEM_IF_CSR_CS_WIDTH: integer := 3
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_rst_n       : in     vl_logic;
        avalon_mm_addr  : in     vl_logic_vector;
        avalon_mm_be    : in     vl_logic_vector;
        avalon_mm_write : in     vl_logic;
        avalon_mm_wdata : in     vl_logic_vector;
        avalon_mm_read  : in     vl_logic;
        avalon_mm_rdata : out    vl_logic_vector;
        avalon_mm_rdata_valid: out    vl_logic;
        avalon_mm_waitrequest: out    vl_logic;
        sts_cal_success : in     vl_logic;
        sts_cal_fail    : in     vl_logic;
        local_power_down_ack: in     vl_logic;
        local_self_rfsh_ack: in     vl_logic;
        sts_sbe_error   : in     vl_logic;
        sts_dbe_error   : in     vl_logic;
        sts_corr_dropped: in     vl_logic;
        sts_sbe_count   : in     vl_logic_vector(7 downto 0);
        sts_dbe_count   : in     vl_logic_vector(7 downto 0);
        sts_corr_dropped_count: in     vl_logic_vector(7 downto 0);
        sts_err_addr    : in     vl_logic_vector(31 downto 0);
        sts_corr_dropped_addr: in     vl_logic_vector(31 downto 0);
        cfg_cal_req     : out    vl_logic;
        cfg_clock_off   : out    vl_logic_vector;
        ctl_cal_byte_lane_sel_n: out    vl_logic_vector;
        cfg_cas_wr_lat  : out    vl_logic_vector;
        cfg_add_lat     : out    vl_logic_vector;
        cfg_tcl         : out    vl_logic_vector;
        cfg_burst_length: out    vl_logic_vector;
        cfg_trrd        : out    vl_logic_vector;
        cfg_tfaw        : out    vl_logic_vector;
        cfg_trfc        : out    vl_logic_vector;
        cfg_trefi       : out    vl_logic_vector;
        cfg_trcd        : out    vl_logic_vector;
        cfg_trp         : out    vl_logic_vector;
        cfg_twr         : out    vl_logic_vector;
        cfg_twtr        : out    vl_logic_vector;
        cfg_trtp        : out    vl_logic_vector;
        cfg_tras        : out    vl_logic_vector;
        cfg_trc         : out    vl_logic_vector;
        cfg_auto_pd_cycles: out    vl_logic_vector;
        cfg_addr_order  : out    vl_logic_vector(1 downto 0);
        cfg_col_addr_width: out    vl_logic_vector;
        cfg_row_addr_width: out    vl_logic_vector;
        cfg_bank_addr_width: out    vl_logic_vector;
        cfg_cs_addr_width: out    vl_logic_vector;
        cfg_enable_ecc  : out    vl_logic;
        cfg_enable_auto_corr: out    vl_logic;
        cfg_gen_sbe     : out    vl_logic;
        cfg_gen_dbe     : out    vl_logic;
        cfg_enable_intr : out    vl_logic;
        cfg_mask_sbe_intr: out    vl_logic;
        cfg_mask_dbe_intr: out    vl_logic;
        cfg_mask_corr_dropped_intr: out    vl_logic;
        cfg_clr_intr    : out    vl_logic;
        cfg_regdimm_enable: out    vl_logic;
        cfg_reorder_data: out    vl_logic;
        cfg_starve_limit: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CTL_CSR_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_CSR_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_CSR_READ_ONLY : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_CSR_READ_ONLY : constant is 1;
    attribute mti_svvh_generic_type of CFG_AVALON_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_AVALON_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CLK_PAIR_COUNT : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of \CFG_CS_ADDR_WIDTH\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_ROW_ADDR_WIDTH\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_COL_ADDR_WIDTH\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_BANK_ADDR_WIDTH\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_ENABLE_ECC\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_ENABLE_AUTO_CORR\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_REGDIMM_ENABLE\ : constant is 1;
    attribute mti_svvh_generic_type of CAS_WR_LAT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ADD_LAT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TCL_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of BL_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRRD_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TFAW_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRFC_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TREFI_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRCD_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRP_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TWR_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TWTR_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRTP_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRAS_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TRC_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AUTO_PD_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of STARVE_LIMIT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of \CFG_CAS_WR_LAT\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_ADD_LAT\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TCL\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_BURST_LENGTH\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRRD\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TFAW\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRFC\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TREFI\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRCD\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRP\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TWR\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TWTR\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRTP\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRAS\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_TRC\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_AUTO_PD_CYCLES\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_ADDR_ORDER\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_REORDER_DATA\ : constant is 1;
    attribute mti_svvh_generic_type of \CFG_STARVE_LIMIT\ : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CSR_COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CSR_ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CSR_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CSR_CS_WIDTH : constant is 1;
end alt_mem_ddrx_csr;
