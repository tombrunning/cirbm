library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_addr_cmd_wrap is
    generic(
        CFG_MEM_IF_CHIP : integer := 2;
        CFG_MEM_IF_CKE_WIDTH: integer := 2;
        CFG_MEM_IF_ADDR_WIDTH: integer := 16;
        CFG_MEM_IF_ROW_WIDTH: integer := 16;
        CFG_MEM_IF_COL_WIDTH: integer := 12;
        CFG_MEM_IF_BA_WIDTH: integer := 3;
        CFG_LPDDR2_ENABLED: integer := 1;
        CFG_PORT_WIDTH_TYPE: integer := 3;
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_AFI_INTF_PHASE_NUM: integer := 2;
        CFG_LOCAL_ID_WIDTH: integer := 8;
        CFG_DATA_ID_WIDTH: integer := 4;
        CFG_INT_SIZE_WIDTH: integer := 4;
        CFG_ODT_ENABLED : integer := 1;
        CFG_MEM_IF_ODT_WIDTH: integer := 2;
        CFG_PORT_WIDTH_CAS_WR_LAT: integer := 5;
        CFG_PORT_WIDTH_TCL: integer := 5;
        CFG_PORT_WIDTH_ADD_LAT: integer := 5;
        CFG_PORT_WIDTH_WRITE_ODT_CHIP: integer := 4;
        CFG_PORT_WIDTH_READ_ODT_CHIP: integer := 4;
        CFG_PORT_WIDTH_OUTPUT_REGD: integer := 2
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        ctl_cal_success : in     vl_logic;
        cfg_type        : in     vl_logic_vector;
        cfg_tcl         : in     vl_logic_vector;
        cfg_cas_wr_lat  : in     vl_logic_vector;
        cfg_add_lat     : in     vl_logic_vector;
        cfg_write_odt_chip: in     vl_logic_vector;
        cfg_read_odt_chip: in     vl_logic_vector;
        cfg_burst_length: in     vl_logic_vector(4 downto 0);
        cfg_output_regd_for_afi_output: in     vl_logic_vector;
        bg_do_write     : in     vl_logic_vector;
        bg_do_read      : in     vl_logic_vector;
        bg_do_burst_chop: in     vl_logic_vector;
        bg_do_burst_terminate: in     vl_logic_vector;
        bg_do_auto_precharge: in     vl_logic_vector;
        bg_do_activate  : in     vl_logic_vector;
        bg_do_precharge : in     vl_logic_vector;
        bg_do_precharge_all: in     vl_logic_vector;
        bg_do_refresh   : in     vl_logic_vector;
        bg_do_self_refresh: in     vl_logic_vector;
        bg_do_power_down: in     vl_logic_vector;
        bg_do_deep_pdown: in     vl_logic_vector;
        bg_do_rmw_correct: in     vl_logic_vector;
        bg_do_rmw_partial: in     vl_logic_vector;
        bg_do_lmr_read  : in     vl_logic;
        bg_do_refresh_1bank: in     vl_logic;
        bg_do_zq_cal    : in     vl_logic_vector;
        bg_do_lmr       : in     vl_logic_vector;
        bg_localid      : in     vl_logic_vector;
        bg_dataid       : in     vl_logic_vector;
        bg_size         : in     vl_logic_vector;
        bg_to_chip      : in     vl_logic_vector;
        bg_to_bank      : in     vl_logic_vector;
        bg_to_row       : in     vl_logic_vector;
        bg_to_col       : in     vl_logic_vector;
        bg_to_lmr       : in     vl_logic_vector(7 downto 0);
        lmr_opcode      : in     vl_logic_vector;
        afi_cke         : out    vl_logic_vector;
        afi_cs_n        : out    vl_logic_vector;
        afi_ras_n       : out    vl_logic_vector;
        afi_cas_n       : out    vl_logic_vector;
        afi_we_n        : out    vl_logic_vector;
        afi_ba          : out    vl_logic_vector;
        afi_addr        : out    vl_logic_vector;
        afi_rst_n       : out    vl_logic_vector;
        afi_odt         : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CKE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_BA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LPDDR2_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_AFI_INTF_PHASE_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_INT_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_ODT_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_CAS_WR_LAT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TCL : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ADD_LAT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_WRITE_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_READ_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_OUTPUT_REGD : constant is 1;
end alt_mem_ddrx_addr_cmd_wrap;
