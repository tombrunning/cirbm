library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_c0 is
    port(
        afi_reset_n     : in     vl_logic;
        afi_clk         : in     vl_logic;
        afi_half_clk    : in     vl_logic;
        local_init_done : out    vl_logic;
        local_cal_success: out    vl_logic;
        local_cal_fail  : out    vl_logic;
        afi_addr        : out    vl_logic_vector(27 downto 0);
        afi_ba          : out    vl_logic_vector(5 downto 0);
        afi_ras_n       : out    vl_logic_vector(1 downto 0);
        afi_we_n        : out    vl_logic_vector(1 downto 0);
        afi_cas_n       : out    vl_logic_vector(1 downto 0);
        afi_odt         : out    vl_logic_vector(1 downto 0);
        afi_cke         : out    vl_logic_vector(1 downto 0);
        afi_cs_n        : out    vl_logic_vector(1 downto 0);
        afi_dqs_burst   : out    vl_logic_vector(15 downto 0);
        afi_wdata_valid : out    vl_logic_vector(15 downto 0);
        afi_wdata       : out    vl_logic_vector(255 downto 0);
        afi_dm          : out    vl_logic_vector(31 downto 0);
        afi_rdata       : in     vl_logic_vector(255 downto 0);
        afi_mem_clk_disable: out    vl_logic_vector(1 downto 0);
        afi_init_req    : out    vl_logic;
        afi_cal_req     : out    vl_logic;
        afi_rdata_en    : out    vl_logic_vector(1 downto 0);
        afi_rdata_en_full: out    vl_logic_vector(1 downto 0);
        afi_rdata_valid : in     vl_logic_vector(1 downto 0);
        afi_cal_success : in     vl_logic;
        afi_cal_fail    : in     vl_logic;
        afi_wlat        : in     vl_logic_vector(5 downto 0);
        afi_rlat        : in     vl_logic_vector(5 downto 0);
        avl_ready       : out    vl_logic;
        avl_burstbegin  : in     vl_logic;
        avl_addr        : in     vl_logic_vector(24 downto 0);
        avl_rdata_valid : out    vl_logic;
        avl_rdata       : out    vl_logic_vector(255 downto 0);
        avl_wdata       : in     vl_logic_vector(255 downto 0);
        avl_be          : in     vl_logic_vector(31 downto 0);
        avl_read_req    : in     vl_logic;
        avl_write_req   : in     vl_logic;
        avl_size        : in     vl_logic_vector(2 downto 0)
    );
end DE4_QSYS_mem_if_ddr2_emif_c0;
