// DE4_QSYS_tb.v

// Generated using ACDS version 13.0sp1 232 at 2015.07.01.13:28:27

`timescale 1 ps / 1 ps
module DE4_QSYS_tb (
	);

	wire         de4_qsys_inst_clk_bfm_clk_clk;                           // DE4_QSYS_inst_clk_bfm:clk -> [DE4_QSYS_inst:clk_clk, DE4_QSYS_inst_reset_bfm:clk]
	wire         de4_qsys_inst_reset_bfm_reset_reset;                     // DE4_QSYS_inst_reset_bfm:reset -> DE4_QSYS_inst:reset_reset_n
	wire         de4_qsys_inst_oct_bfm_conduit_rdn;                       // DE4_QSYS_inst_oct_bfm:sig_rdn -> DE4_QSYS_inst:oct_rdn
	wire         de4_qsys_inst_oct_bfm_conduit_rup;                       // DE4_QSYS_inst_oct_bfm:sig_rup -> DE4_QSYS_inst:oct_rup
	wire         de4_qsys_inst_mem_if_ddr2_emif_status_local_cal_fail;    // DE4_QSYS_inst:mem_if_ddr2_emif_status_local_cal_fail -> DE4_QSYS_inst_mem_if_ddr2_emif_status_bfm:sig_local_cal_fail
	wire         de4_qsys_inst_mem_if_ddr2_emif_status_local_cal_success; // DE4_QSYS_inst:mem_if_ddr2_emif_status_local_cal_success -> DE4_QSYS_inst_mem_if_ddr2_emif_status_bfm:sig_local_cal_success
	wire         de4_qsys_inst_mem_if_ddr2_emif_status_local_init_done;   // DE4_QSYS_inst:mem_if_ddr2_emif_status_local_init_done -> DE4_QSYS_inst_mem_if_ddr2_emif_status_bfm:sig_local_init_done
	wire   [7:0] de4_qsys_inst_led_export;                                // DE4_QSYS_inst:led_export -> DE4_QSYS_inst_led_bfm:sig_export
	wire   [3:0] de4_qsys_inst_button_bfm_conduit_export;                 // DE4_QSYS_inst_button_bfm:sig_export -> DE4_QSYS_inst:button_export
	wire         de4_qsys_inst_ddr2_i2c_scl_export;                       // DE4_QSYS_inst:ddr2_i2c_scl_export -> DE4_QSYS_inst_ddr2_i2c_scl_bfm:sig_export
	wire         de4_qsys_inst_ddr2_i2c_sda_export;                       // [] -> [DE4_QSYS_inst:ddr2_i2c_sda_export, DE4_QSYS_inst_ddr2_i2c_sda_bfm:sig_export]
	wire   [0:0] de4_qsys_inst_memory_mem_odt;                            // DE4_QSYS_inst:memory_mem_odt -> mem_if_ddr2_emif_mem_model:mem_odt
	wire   [0:0] de4_qsys_inst_memory_mem_cs_n;                           // DE4_QSYS_inst:memory_mem_cs_n -> mem_if_ddr2_emif_mem_model:mem_cs_n
	wire  [13:0] de4_qsys_inst_memory_mem_a;                              // DE4_QSYS_inst:memory_mem_a -> mem_if_ddr2_emif_mem_model:mem_a
	wire   [1:0] de4_qsys_inst_memory_mem_ck_n;                           // DE4_QSYS_inst:memory_mem_ck_n -> mem_if_ddr2_emif_mem_model:mem_ck_n
	wire   [0:0] de4_qsys_inst_memory_mem_ras_n;                          // DE4_QSYS_inst:memory_mem_ras_n -> mem_if_ddr2_emif_mem_model:mem_ras_n
	wire   [0:0] de4_qsys_inst_memory_mem_cke;                            // DE4_QSYS_inst:memory_mem_cke -> mem_if_ddr2_emif_mem_model:mem_cke
	wire   [7:0] de4_qsys_inst_memory_mem_dqs;                            // [] -> [DE4_QSYS_inst:memory_mem_dqs, mem_if_ddr2_emif_mem_model:mem_dqs]
	wire   [0:0] de4_qsys_inst_memory_mem_we_n;                           // DE4_QSYS_inst:memory_mem_we_n -> mem_if_ddr2_emif_mem_model:mem_we_n
	wire   [2:0] de4_qsys_inst_memory_mem_ba;                             // DE4_QSYS_inst:memory_mem_ba -> mem_if_ddr2_emif_mem_model:mem_ba
	wire  [63:0] de4_qsys_inst_memory_mem_dq;                             // [] -> [DE4_QSYS_inst:memory_mem_dq, mem_if_ddr2_emif_mem_model:mem_dq]
	wire   [1:0] de4_qsys_inst_memory_mem_ck;                             // DE4_QSYS_inst:memory_mem_ck -> mem_if_ddr2_emif_mem_model:mem_ck
	wire   [7:0] de4_qsys_inst_memory_mem_dm;                             // DE4_QSYS_inst:memory_mem_dm -> mem_if_ddr2_emif_mem_model:mem_dm
	wire   [0:0] de4_qsys_inst_memory_mem_cas_n;                          // DE4_QSYS_inst:memory_mem_cas_n -> mem_if_ddr2_emif_mem_model:mem_cas_n
	wire   [7:0] de4_qsys_inst_memory_mem_dqs_n;                          // [] -> [DE4_QSYS_inst:memory_mem_dqs_n, mem_if_ddr2_emif_mem_model:mem_dqs_n]

	DE4_QSYS de4_qsys_inst (
		.clk_clk                                   (de4_qsys_inst_clk_bfm_clk_clk),                           //                     clk.clk
		.reset_reset_n                             (de4_qsys_inst_reset_bfm_reset_reset),                     //                   reset.reset_n
		.memory_mem_a                              (de4_qsys_inst_memory_mem_a),                              //                  memory.mem_a
		.memory_mem_ba                             (de4_qsys_inst_memory_mem_ba),                             //                        .mem_ba
		.memory_mem_ck                             (de4_qsys_inst_memory_mem_ck),                             //                        .mem_ck
		.memory_mem_ck_n                           (de4_qsys_inst_memory_mem_ck_n),                           //                        .mem_ck_n
		.memory_mem_cke                            (de4_qsys_inst_memory_mem_cke),                            //                        .mem_cke
		.memory_mem_cs_n                           (de4_qsys_inst_memory_mem_cs_n),                           //                        .mem_cs_n
		.memory_mem_dm                             (de4_qsys_inst_memory_mem_dm),                             //                        .mem_dm
		.memory_mem_ras_n                          (de4_qsys_inst_memory_mem_ras_n),                          //                        .mem_ras_n
		.memory_mem_cas_n                          (de4_qsys_inst_memory_mem_cas_n),                          //                        .mem_cas_n
		.memory_mem_we_n                           (de4_qsys_inst_memory_mem_we_n),                           //                        .mem_we_n
		.memory_mem_dq                             (de4_qsys_inst_memory_mem_dq),                             //                        .mem_dq
		.memory_mem_dqs                            (de4_qsys_inst_memory_mem_dqs),                            //                        .mem_dqs
		.memory_mem_dqs_n                          (de4_qsys_inst_memory_mem_dqs_n),                          //                        .mem_dqs_n
		.memory_mem_odt                            (de4_qsys_inst_memory_mem_odt),                            //                        .mem_odt
		.oct_rdn                                   (de4_qsys_inst_oct_bfm_conduit_rdn),                       //                     oct.rdn
		.oct_rup                                   (de4_qsys_inst_oct_bfm_conduit_rup),                       //                        .rup
		.mem_if_ddr2_emif_status_local_init_done   (de4_qsys_inst_mem_if_ddr2_emif_status_local_init_done),   // mem_if_ddr2_emif_status.local_init_done
		.mem_if_ddr2_emif_status_local_cal_success (de4_qsys_inst_mem_if_ddr2_emif_status_local_cal_success), //                        .local_cal_success
		.mem_if_ddr2_emif_status_local_cal_fail    (de4_qsys_inst_mem_if_ddr2_emif_status_local_cal_fail),    //                        .local_cal_fail
		.led_export                                (de4_qsys_inst_led_export),                                //                     led.export
		.button_export                             (de4_qsys_inst_button_bfm_conduit_export),                 //                  button.export
		.ddr2_i2c_scl_export                       (de4_qsys_inst_ddr2_i2c_scl_export),                       //            ddr2_i2c_scl.export
		.ddr2_i2c_sda_export                       (de4_qsys_inst_ddr2_i2c_sda_export)                        //            ddr2_i2c_sda.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) de4_qsys_inst_clk_bfm (
		.clk (de4_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) de4_qsys_inst_reset_bfm (
		.reset (de4_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (de4_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm de4_qsys_inst_oct_bfm (
		.sig_rdn (de4_qsys_inst_oct_bfm_conduit_rdn), // conduit.rdn
		.sig_rup (de4_qsys_inst_oct_bfm_conduit_rup)  //        .rup
	);

	altera_conduit_bfm_0002 de4_qsys_inst_mem_if_ddr2_emif_status_bfm (
		.sig_local_init_done   (de4_qsys_inst_mem_if_ddr2_emif_status_local_init_done),   // conduit.local_init_done
		.sig_local_cal_success (de4_qsys_inst_mem_if_ddr2_emif_status_local_cal_success), //        .local_cal_success
		.sig_local_cal_fail    (de4_qsys_inst_mem_if_ddr2_emif_status_local_cal_fail)     //        .local_cal_fail
	);

	altera_conduit_bfm_0003 de4_qsys_inst_led_bfm (
		.sig_export (de4_qsys_inst_led_export)  // conduit.export
	);

	altera_conduit_bfm_0004 de4_qsys_inst_button_bfm (
		.sig_export (de4_qsys_inst_button_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0005 de4_qsys_inst_ddr2_i2c_scl_bfm (
		.sig_export (de4_qsys_inst_ddr2_i2c_scl_export)  // conduit.export
	);

	altera_conduit_bfm_0006 de4_qsys_inst_ddr2_i2c_sda_bfm (
		.sig_export (de4_qsys_inst_ddr2_i2c_sda_export)  // conduit.export
	);

	alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en #(
		.MEM_IF_ADDR_WIDTH            (14),
		.MEM_IF_ROW_ADDR_WIDTH        (14),
		.MEM_IF_COL_ADDR_WIDTH        (10),
		.MEM_IF_CS_PER_RANK           (1),
		.MEM_IF_CONTROL_WIDTH         (1),
		.MEM_IF_DQS_WIDTH             (8),
		.MEM_IF_CS_WIDTH              (1),
		.MEM_IF_BANKADDR_WIDTH        (3),
		.MEM_IF_DQ_WIDTH              (64),
		.MEM_IF_CK_WIDTH              (2),
		.MEM_IF_CLK_EN_WIDTH          (1),
		.DEVICE_WIDTH                 (1),
		.MEM_TRCD                     (5),
		.MEM_TRTP                     (3),
		.MEM_DQS_TO_CLK_CAPTURE_DELAY (100),
		.MEM_CLK_TO_DQS_CAPTURE_DELAY (100000),
		.MEM_IF_ODT_WIDTH             (1),
		.MEM_MIRROR_ADDRESSING_DEC    (0),
		.MEM_REGDIMM_ENABLED          (0),
		.DEVICE_DEPTH                 (1),
		.MEM_GUARANTEED_WRITE_INIT    (0),
		.MEM_VERBOSE                  (1),
		.MEM_INIT_EN                  (0),
		.MEM_INIT_FILE                (""),
		.DAT_DATA_WIDTH               (32)
	) mem_if_ddr2_emif_mem_model (
		.mem_a     (de4_qsys_inst_memory_mem_a),     // memory.mem_a
		.mem_ba    (de4_qsys_inst_memory_mem_ba),    //       .mem_ba
		.mem_ck    (de4_qsys_inst_memory_mem_ck),    //       .mem_ck
		.mem_ck_n  (de4_qsys_inst_memory_mem_ck_n),  //       .mem_ck_n
		.mem_cke   (de4_qsys_inst_memory_mem_cke),   //       .mem_cke
		.mem_cs_n  (de4_qsys_inst_memory_mem_cs_n),  //       .mem_cs_n
		.mem_dm    (de4_qsys_inst_memory_mem_dm),    //       .mem_dm
		.mem_ras_n (de4_qsys_inst_memory_mem_ras_n), //       .mem_ras_n
		.mem_cas_n (de4_qsys_inst_memory_mem_cas_n), //       .mem_cas_n
		.mem_we_n  (de4_qsys_inst_memory_mem_we_n),  //       .mem_we_n
		.mem_dq    (de4_qsys_inst_memory_mem_dq),    //       .mem_dq
		.mem_dqs   (de4_qsys_inst_memory_mem_dqs),   //       .mem_dqs
		.mem_dqs_n (de4_qsys_inst_memory_mem_dqs_n), //       .mem_dqs_n
		.mem_odt   (de4_qsys_inst_memory_mem_odt)    //       .mem_odt
	);

endmodule
