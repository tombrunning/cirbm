library verilog;
use verilog.vl_types.all;
entity altera_conduit_bfm_0003 is
    port(
        sig_export      : in     vl_logic_vector(7 downto 0)
    );
end altera_conduit_bfm_0003;
