library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_pll0 is
    generic(
        DEVICE_FAMILY   : string  := "Stratix IV";
        ALTERA_ALT_MEM_IF_PHY_FAST_SIM_MODEL: integer := 1;
        PLL_PHASE_COUNTER_WIDTH: integer := 4;
        GENERIC_PLL     : string  := "false";
        REF_CLK_FREQ    : string  := "50.0 MHz";
        REF_CLK_PERIOD_PS: integer := 20000;
        PLL_AFI_CLK_FREQ_STR: string  := "150.0 MHz";
        PLL_MEM_CLK_FREQ_STR: string  := "300.0 MHz";
        PLL_WRITE_CLK_FREQ_STR: string  := "300.0 MHz";
        PLL_ADDR_CMD_CLK_FREQ_STR: string  := "150.0 MHz";
        PLL_AFI_HALF_CLK_FREQ_STR: string  := "75.0 MHz";
        PLL_NIOS_CLK_FREQ_STR: string  := "75.0 MHz";
        PLL_CONFIG_CLK_FREQ_STR: string  := "25.0 MHz";
        PLL_P2C_READ_CLK_FREQ_STR: string  := "";
        PLL_C2P_WRITE_CLK_FREQ_STR: string  := "";
        PLL_HR_CLK_FREQ_STR: string  := "";
        PLL_DR_CLK_FREQ_STR: string  := "";
        PLL_AFI_CLK_FREQ_SIM_STR: string  := "6668 ps";
        PLL_MEM_CLK_FREQ_SIM_STR: string  := "3334 ps";
        PLL_WRITE_CLK_FREQ_SIM_STR: string  := "3334 ps";
        PLL_ADDR_CMD_CLK_FREQ_SIM_STR: string  := "6668 ps";
        PLL_AFI_HALF_CLK_FREQ_SIM_STR: string  := "13336 ps";
        PLL_NIOS_CLK_FREQ_SIM_STR: string  := "13336 ps";
        PLL_CONFIG_CLK_FREQ_SIM_STR: string  := "40008 ps";
        PLL_P2C_READ_CLK_FREQ_SIM_STR: string  := "0 ps";
        PLL_C2P_WRITE_CLK_FREQ_SIM_STR: string  := "0 ps";
        PLL_HR_CLK_FREQ_SIM_STR: string  := "0 ps";
        PLL_DR_CLK_FREQ_SIM_STR: string  := "0 ps";
        AFI_CLK_PHASE   : string  := "0 ps";
        MEM_CLK_PHASE   : string  := "0 ps";
        WRITE_CLK_PHASE : string  := "833 ps";
        ADDR_CMD_CLK_PHASE: string  := "5000 ps";
        AFI_HALF_CLK_PHASE: string  := "0 ps";
        AVL_CLK_PHASE   : string  := "0 ps";
        CONFIG_CLK_PHASE: string  := "0 ps";
        ABSTRACT_REAL_COMPARE_TEST: string  := "false";
        PLL_AFI_CLK_DIV : integer := 1;
        PLL_MEM_CLK_DIV : integer := 1;
        PLL_WRITE_CLK_DIV: integer := 1;
        PLL_ADDR_CMD_CLK_DIV: integer := 1;
        PLL_AFI_HALF_CLK_DIV: integer := 2;
        PLL_NIOS_CLK_DIV: integer := 2;
        PLL_CONFIG_CLK_DIV: integer := 2;
        PLL_AFI_CLK_MULT: integer := 3;
        PLL_MEM_CLK_MULT: integer := 6;
        PLL_WRITE_CLK_MULT: integer := 6;
        PLL_ADDR_CMD_CLK_MULT: integer := 3;
        PLL_AFI_HALF_CLK_MULT: integer := 3;
        PLL_NIOS_CLK_MULT: integer := 3;
        PLL_CONFIG_CLK_MULT: integer := 1;
        PLL_AFI_CLK_PHASE_PS: string  := "0";
        PLL_MEM_CLK_PHASE_PS: string  := "0";
        PLL_WRITE_CLK_PHASE_PS: string  := "833";
        PLL_ADDR_CMD_CLK_PHASE_PS: string  := "5000";
        PLL_AFI_HALF_CLK_PHASE_PS: string  := "0";
        PLL_NIOS_CLK_PHASE_PS: string  := "0";
        PLL_CONFIG_CLK_PHASE_PS: string  := "0"
    );
    port(
        global_reset_n  : in     vl_logic;
        pll_ref_clk     : in     vl_logic;
        pll_mem_clk     : out    vl_logic;
        pll_write_clk   : out    vl_logic;
        pll_write_clk_pre_phy_clk: out    vl_logic;
        pll_addr_cmd_clk: out    vl_logic;
        pll_avl_clk     : out    vl_logic;
        pll_config_clk  : out    vl_logic;
        pll_locked      : out    vl_logic;
        afi_clk         : out    vl_logic;
        afi_half_clk    : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of ALTERA_ALT_MEM_IF_PHY_FAST_SIM_MODEL : constant is 1;
    attribute mti_svvh_generic_type of PLL_PHASE_COUNTER_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of GENERIC_PLL : constant is 1;
    attribute mti_svvh_generic_type of REF_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of REF_CLK_PERIOD_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_MEM_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_WRITE_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_ADDR_CMD_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_HALF_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_NIOS_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_CONFIG_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_P2C_READ_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_C2P_WRITE_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_HR_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_DR_CLK_FREQ_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_MEM_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_WRITE_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_ADDR_CMD_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_HALF_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_NIOS_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_CONFIG_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_P2C_READ_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_C2P_WRITE_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_HR_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of PLL_DR_CLK_FREQ_SIM_STR : constant is 1;
    attribute mti_svvh_generic_type of AFI_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of WRITE_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of ADDR_CMD_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of AFI_HALF_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of AVL_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of CONFIG_CLK_PHASE : constant is 1;
    attribute mti_svvh_generic_type of ABSTRACT_REAL_COMPARE_TEST : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_MEM_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_WRITE_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_ADDR_CMD_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_HALF_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_NIOS_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_CONFIG_CLK_DIV : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_MEM_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_WRITE_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_ADDR_CMD_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_HALF_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_NIOS_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_CONFIG_CLK_MULT : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_CLK_PHASE_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_MEM_CLK_PHASE_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_WRITE_CLK_PHASE_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_ADDR_CMD_CLK_PHASE_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_AFI_HALF_CLK_PHASE_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_NIOS_CLK_PHASE_PS : constant is 1;
    attribute mti_svvh_generic_type of PLL_CONFIG_CLK_PHASE_PS : constant is 1;
end DE4_QSYS_mem_if_ddr2_emif_pll0;
