library verilog;
use verilog.vl_types.all;
entity afi_mux_ddrx is
    generic(
        AFI_ADDR_WIDTH  : integer := 0;
        AFI_BANKADDR_WIDTH: integer := 0;
        AFI_CS_WIDTH    : integer := 0;
        AFI_CLK_EN_WIDTH: integer := 0;
        AFI_ODT_WIDTH   : integer := 0;
        AFI_WLAT_WIDTH  : integer := 0;
        AFI_RLAT_WIDTH  : integer := 0;
        AFI_DM_WIDTH    : integer := 0;
        AFI_CONTROL_WIDTH: integer := 0;
        AFI_DQ_WIDTH    : integer := 0;
        AFI_WRITE_DQS_WIDTH: integer := 0;
        AFI_RATE_RATIO  : integer := 0;
        MRS_MIRROR_PING_PONG_ATSO: integer := 0
    );
    port(
        clk             : in     vl_logic;
        mux_sel         : in     vl_logic;
        afi_addr        : in     vl_logic_vector;
        afi_ba          : in     vl_logic_vector;
        afi_cs_n        : in     vl_logic_vector;
        afi_cke         : in     vl_logic_vector;
        afi_odt         : in     vl_logic_vector;
        afi_ras_n       : in     vl_logic_vector;
        afi_cas_n       : in     vl_logic_vector;
        afi_we_n        : in     vl_logic_vector;
        afi_dm          : in     vl_logic_vector;
        afi_wlat        : out    vl_logic_vector;
        afi_rlat        : out    vl_logic_vector;
        afi_dqs_burst   : in     vl_logic_vector;
        afi_wdata       : in     vl_logic_vector;
        afi_wdata_valid : in     vl_logic_vector;
        afi_rdata_en    : in     vl_logic_vector;
        afi_rdata_en_full: in     vl_logic_vector;
        afi_rdata       : out    vl_logic_vector;
        afi_rdata_valid : out    vl_logic_vector;
        afi_cal_success : out    vl_logic;
        afi_cal_fail    : out    vl_logic;
        seq_mux_addr    : in     vl_logic_vector;
        seq_mux_ba      : in     vl_logic_vector;
        seq_mux_cs_n    : in     vl_logic_vector;
        seq_mux_cke     : in     vl_logic_vector;
        seq_mux_odt     : in     vl_logic_vector;
        seq_mux_ras_n   : in     vl_logic_vector;
        seq_mux_cas_n   : in     vl_logic_vector;
        seq_mux_we_n    : in     vl_logic_vector;
        seq_mux_dm      : in     vl_logic_vector;
        seq_mux_dqs_burst: in     vl_logic_vector;
        seq_mux_wdata   : in     vl_logic_vector;
        seq_mux_wdata_valid: in     vl_logic_vector;
        seq_mux_rdata_en: in     vl_logic_vector;
        seq_mux_rdata_en_full: in     vl_logic_vector;
        seq_mux_rdata   : out    vl_logic_vector;
        seq_mux_rdata_valid: out    vl_logic_vector;
        phy_mux_addr    : out    vl_logic_vector;
        phy_mux_ba      : out    vl_logic_vector;
        phy_mux_cs_n    : out    vl_logic_vector;
        phy_mux_cke     : out    vl_logic_vector;
        phy_mux_odt     : out    vl_logic_vector;
        phy_mux_ras_n   : out    vl_logic_vector;
        phy_mux_cas_n   : out    vl_logic_vector;
        phy_mux_we_n    : out    vl_logic_vector;
        phy_mux_dm      : out    vl_logic_vector;
        phy_mux_wlat    : in     vl_logic_vector;
        phy_mux_rlat    : in     vl_logic_vector;
        phy_mux_dqs_burst: out    vl_logic_vector;
        phy_mux_wdata   : out    vl_logic_vector;
        phy_mux_wdata_valid: out    vl_logic_vector;
        phy_mux_rdata_en: out    vl_logic_vector;
        phy_mux_rdata_en_full: out    vl_logic_vector;
        phy_mux_rdata   : in     vl_logic_vector;
        phy_mux_rdata_valid: in     vl_logic_vector;
        phy_mux_cal_success: in     vl_logic;
        phy_mux_cal_fail: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AFI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_WLAT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RLAT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATE_RATIO : constant is 1;
    attribute mti_svvh_generic_type of MRS_MIRROR_PING_PONG_ATSO : constant is 1;
end afi_mux_ddrx;
