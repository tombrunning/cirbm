library verilog;
use verilog.vl_types.all;
entity mem_rank_model is
    generic(
        MEM_IF_BA_WIDTH : integer := 2;
        MEM_IF_ADDR_WIDTH: integer := 12;
        MEM_IF_ROW_ADDR_WIDTH: integer := 12;
        MEM_IF_COL_ADDR_WIDTH: integer := 10;
        MEM_DQS_WIDTH   : integer := 2;
        MEM_DQ_WIDTH    : integer := 16;
        MEM_TRTP        : integer := 6;
        MEM_TRCD        : integer := 11;
        MEM_DQS_TO_CLK_CAPTURE_DELAY: integer := 0;
        MEM_CLK_TO_DQS_CAPTURE_DELAY: integer := 0;
        MEM_MIRROR_ADDRESSING: integer := 0;
        MEM_DEPTH_IDX   : integer := -1;
        MEM_WIDTH_IDX   : integer := -1;
        MEM_RANK_IDX    : integer := -1;
        MEM_INIT_EN     : integer := 0;
        MEM_INIT_FILE   : string  := "";
        MEM_GUARANTEED_WRITE_INIT: integer := 0;
        DAT_DATA_WIDTH  : integer := 32;
        MEM_VERBOSE     : integer := 1;
        REFRESH_BURST_VALIDATION: integer := 0
    );
    port(
        mem_a           : in     vl_logic_vector;
        mem_ba          : in     vl_logic_vector;
        mem_ck          : in     vl_logic;
        mem_ck_n        : in     vl_logic;
        mem_cke         : in     vl_logic;
        mem_ras_n       : in     vl_logic;
        mem_cas_n       : in     vl_logic;
        mem_we_n        : in     vl_logic;
        mem_dm          : in     vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        mem_odt         : in     vl_logic;
        mem_cs_n        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MEM_IF_BA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ROW_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_COL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRTP : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRCD : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_TO_CLK_CAPTURE_DELAY : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_TO_DQS_CAPTURE_DELAY : constant is 1;
    attribute mti_svvh_generic_type of MEM_MIRROR_ADDRESSING : constant is 1;
    attribute mti_svvh_generic_type of MEM_DEPTH_IDX : constant is 1;
    attribute mti_svvh_generic_type of MEM_WIDTH_IDX : constant is 1;
    attribute mti_svvh_generic_type of MEM_RANK_IDX : constant is 1;
    attribute mti_svvh_generic_type of MEM_INIT_EN : constant is 1;
    attribute mti_svvh_generic_type of MEM_INIT_FILE : constant is 1;
    attribute mti_svvh_generic_type of MEM_GUARANTEED_WRITE_INIT : constant is 1;
    attribute mti_svvh_generic_type of DAT_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_VERBOSE : constant is 1;
    attribute mti_svvh_generic_type of REFRESH_BURST_VALIDATION : constant is 1;
end mem_rank_model;
