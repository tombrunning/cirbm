library verilog;
use verilog.vl_types.all;
entity alt_mem_if_nextgen_ddr2_controller_core is
    generic(
        AVL_SIZE_WIDTH  : integer := 0;
        AVL_ADDR_WIDTH  : integer := 0;
        AVL_DATA_WIDTH  : integer := 0;
        LOCAL_ID_WIDTH  : integer := 0;
        AVL_BE_WIDTH    : integer := 0;
        LOCAL_CS_WIDTH  : integer := 0;
        MEM_IF_ADDR_WIDTH: integer := 0;
        MEM_IF_CLK_PAIR_COUNT: integer := 0;
        LOCAL_IF_TYPE   : string  := "AVALON";
        DWIDTH_RATIO    : integer := 0;
        CTL_ODT_ENABLED : integer := 0;
        CTL_OUTPUT_REGD : integer := 0;
        CTL_TBP_NUM     : integer := 0;
        WRBUFFER_ADDR_WIDTH: integer := 0;
        RDBUFFER_ADDR_WIDTH: integer := 0;
        MEM_IF_CS_WIDTH : integer := 0;
        MEM_IF_CHIP_BITS: integer := 0;
        MEM_IF_BANKADDR_WIDTH: integer := 0;
        MEM_IF_ROW_ADDR_WIDTH: integer := 0;
        MEM_IF_COL_ADDR_WIDTH: integer := 0;
        MEM_IF_ODT_WIDTH: integer := 0;
        MEM_IF_CLK_EN_WIDTH: integer := 0;
        MEM_IF_DQS_WIDTH: integer := 0;
        MEM_IF_DQ_WIDTH : integer := 0;
        MEM_IF_DM_WIDTH : integer := 0;
        MAX_MEM_IF_CS_WIDTH: integer := 30;
        MAX_MEM_IF_CHIP : integer := 4;
        MAX_MEM_IF_BANKADDR_WIDTH: integer := 3;
        MAX_MEM_IF_ROWADDR_WIDTH: integer := 16;
        MAX_MEM_IF_COLADDR_WIDTH: integer := 12;
        MAX_MEM_IF_ODT_WIDTH: integer := 1;
        MAX_MEM_IF_DQS_WIDTH: integer := 5;
        MAX_MEM_IF_DQ_WIDTH: integer := 40;
        MAX_MEM_IF_MASK_WIDTH: integer := 5;
        MAX_LOCAL_DATA_WIDTH: integer := 80;
        CFG_TYPE        : integer := 0;
        CFG_INTERFACE_WIDTH: integer := 0;
        CFG_BURST_LENGTH: integer := 0;
        CFG_REORDER_DATA: integer := 0;
        CFG_DATA_REORDERING_TYPE: string  := "INTER_ROW";
        CFG_STARVE_LIMIT: integer := 0;
        CFG_ADDR_ORDER  : integer := 0;
        MEM_WTCL_INT    : integer := 0;
        MEM_ADD_LAT     : integer := 0;
        MEM_TCL         : integer := 0;
        MEM_TRRD        : integer := 0;
        MEM_TFAW        : integer := 0;
        MEM_TRFC        : integer := 0;
        MEM_TREFI       : integer := 0;
        MEM_TRCD        : integer := 0;
        MEM_TRP         : integer := 0;
        MEM_TWR         : integer := 0;
        MEM_TWTR        : integer := 0;
        MEM_TRTP        : integer := 0;
        MEM_TRAS        : integer := 0;
        MEM_TRC         : integer := 0;
        CFG_TCCD        : integer := 2;
        MEM_AUTO_PD_CYCLES: integer := 0;
        MEM_IF_RD_TO_WR_TURNAROUND_OCT: integer := 0;
        MEM_IF_WR_TO_RD_TURNAROUND_OCT: integer := 0;
        CTL_RD_TO_PCH_EXTRA_CLK: integer := 0;
        CTL_RD_TO_RD_DIFF_CHIP_EXTRA_CLK: integer := 0;
        CTL_WR_TO_WR_DIFF_CHIP_EXTRA_CLK: integer := 0;
        AFI_ADDR_WIDTH  : integer := 0;
        AFI_BANKADDR_WIDTH: integer := 0;
        AFI_CONTROL_WIDTH: integer := 0;
        AFI_CS_WIDTH    : integer := 0;
        AFI_CLK_EN_WIDTH: integer := 0;
        AFI_ODT_WIDTH   : integer := 0;
        AFI_DM_WIDTH    : integer := 0;
        AFI_DQ_WIDTH    : integer := 0;
        AFI_WRITE_DQS_WIDTH: integer := 0;
        AFI_RATE_RATIO  : integer := 0;
        AFI_WLAT_WIDTH  : integer := 0;
        AFI_RLAT_WIDTH  : integer := 0;
        AFI_RRANK_WIDTH : integer := 0;
        AFI_WRANK_WIDTH : integer := 0;
        USE_SHADOW_REGS : integer := 0;
        CFG_SELF_RFSH_EXIT_CYCLES: integer := 0;
        CFG_PDN_EXIT_CYCLES: integer := 0;
        CFG_POWER_SAVING_EXIT_CYCLES: integer := 0;
        CFG_MEM_CLK_ENTRY_CYCLES: integer := 0;
        MEM_TMRD_CK     : integer := 0;
        CTL_ECC_ENABLED : integer := 0;
        CTL_ECC_AUTO_CORRECTION_ENABLED: integer := 0;
        CTL_ECC_MULTIPLES_16_24_40_72: integer := 1;
        CTL_ENABLE_BURST_INTERRUPT_INT: integer := 0;
        CTL_ENABLE_BURST_TERMINATE_INT: integer := 0;
        CTL_ENABLE_WDATA_PATH_LATENCY: integer := 0;
        CFG_GEN_SBE     : integer := 0;
        CFG_GEN_DBE     : integer := 0;
        CFG_ENABLE_INTR : integer := 0;
        CFG_MASK_SBE_INTR: integer := 0;
        CFG_MASK_DBE_INTR: integer := 0;
        CFG_MASK_CORRDROP_INTR: integer := 0;
        CFG_CLR_INTR    : integer := 0;
        CTL_USR_REFRESH : integer := 0;
        CTL_REGDIMM_ENABLED: integer := 0;
        CFG_WRITE_ODT_CHIP: integer := 0;
        CFG_READ_ODT_CHIP: integer := 0;
        CFG_PORT_WIDTH_WRITE_ODT_CHIP: integer := 0;
        CFG_PORT_WIDTH_READ_ODT_CHIP: integer := 0;
        MEM_IF_CKE_WIDTH: integer := 0;
        CFG_ENABLE_NO_DM: integer := 0;
        CSR_BE_WIDTH    : integer := 4;
        CFG_ERRCMD_FIFO_REG: integer := 0;
        CFG_ECC_DECODER_REG: integer := 0;
        CTL_CSR_ENABLED : integer := 0;
        CSR_ADDR_WIDTH  : integer := 8;
        CSR_DATA_WIDTH  : integer := 32;
        ENABLE_BURST_MERGE: integer := 0
    );
    port(
        afi_clk         : in     vl_logic;
        afi_reset_n     : in     vl_logic;
        afi_half_clk    : in     vl_logic;
        itf_cmd_ready   : out    vl_logic;
        itf_cmd_valid   : in     vl_logic;
        itf_cmd         : in     vl_logic;
        itf_cmd_address : in     vl_logic_vector;
        itf_cmd_burstlen: in     vl_logic_vector;
        itf_cmd_id      : in     vl_logic_vector;
        itf_cmd_priority: in     vl_logic;
        itf_cmd_autopercharge: in     vl_logic;
        itf_cmd_multicast: in     vl_logic;
        itf_wr_data_ready: out    vl_logic;
        itf_wr_data_valid: in     vl_logic;
        itf_wr_data     : in     vl_logic_vector;
        itf_wr_data_byte_en: in     vl_logic_vector;
        itf_wr_data_begin: in     vl_logic;
        itf_wr_data_last: in     vl_logic;
        itf_wr_data_id  : in     vl_logic_vector;
        itf_rd_data_ready: in     vl_logic;
        itf_rd_data_valid: out    vl_logic;
        itf_rd_data     : out    vl_logic_vector;
        itf_rd_data_error: out    vl_logic;
        itf_rd_data_begin: out    vl_logic;
        itf_rd_data_last: out    vl_logic;
        itf_rd_data_id  : out    vl_logic_vector;
        afi_cs_n        : out    vl_logic_vector;
        afi_cke         : out    vl_logic_vector;
        afi_odt         : out    vl_logic_vector;
        afi_addr        : out    vl_logic_vector;
        afi_ba          : out    vl_logic_vector;
        afi_ras_n       : out    vl_logic_vector;
        afi_cas_n       : out    vl_logic_vector;
        afi_we_n        : out    vl_logic_vector;
        afi_dqs_burst   : out    vl_logic_vector;
        afi_wdata_valid : out    vl_logic_vector;
        afi_wdata       : out    vl_logic_vector;
        afi_dm          : out    vl_logic_vector;
        afi_wlat        : in     vl_logic_vector;
        afi_rdata_en    : out    vl_logic_vector;
        afi_rdata_en_full: out    vl_logic_vector;
        afi_rdata       : in     vl_logic_vector;
        afi_rdata_valid : in     vl_logic_vector;
        afi_rlat        : in     vl_logic_vector;
        afi_cal_success : in     vl_logic;
        afi_cal_fail    : in     vl_logic;
        afi_cal_req     : out    vl_logic;
        afi_init_req    : out    vl_logic;
        afi_mem_clk_disable: out    vl_logic_vector;
        local_refresh_ack: out    vl_logic;
        local_powerdn_ack: out    vl_logic;
        local_self_rfsh_ack: out    vl_logic;
        local_deep_powerdn_ack: out    vl_logic;
        local_refresh_req: in     vl_logic;
        local_refresh_chip: in     vl_logic_vector;
        local_self_rfsh_req: in     vl_logic;
        local_self_rfsh_chip: in     vl_logic_vector;
        local_deep_powerdn_req: in     vl_logic;
        local_deep_powerdn_chip: in     vl_logic_vector;
        local_multicast : in     vl_logic;
        local_priority  : in     vl_logic;
        local_init_done : out    vl_logic;
        local_cal_success: out    vl_logic;
        local_cal_fail  : out    vl_logic;
        ecc_interrupt   : out    vl_logic;
        csr_read_req    : in     vl_logic;
        csr_write_req   : in     vl_logic;
        csr_addr        : in     vl_logic_vector;
        csr_wdata       : in     vl_logic_vector;
        csr_rdata       : out    vl_logic_vector;
        csr_be          : in     vl_logic_vector;
        csr_rdata_valid : out    vl_logic;
        csr_waitrequest : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AVL_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AVL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AVL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AVL_BE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CLK_PAIR_COUNT : constant is 1;
    attribute mti_svvh_generic_type of LOCAL_IF_TYPE : constant is 1;
    attribute mti_svvh_generic_type of DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CTL_ODT_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_OUTPUT_REGD : constant is 1;
    attribute mti_svvh_generic_type of CTL_TBP_NUM : constant is 1;
    attribute mti_svvh_generic_type of WRBUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of RDBUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CHIP_BITS : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ROW_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_COL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_ROWADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_COLADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_MEM_IF_MASK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_INTERFACE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_BURST_LENGTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_REORDER_DATA : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_REORDERING_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_STARVE_LIMIT : constant is 1;
    attribute mti_svvh_generic_type of CFG_ADDR_ORDER : constant is 1;
    attribute mti_svvh_generic_type of MEM_WTCL_INT : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADD_LAT : constant is 1;
    attribute mti_svvh_generic_type of MEM_TCL : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRRD : constant is 1;
    attribute mti_svvh_generic_type of MEM_TFAW : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRFC : constant is 1;
    attribute mti_svvh_generic_type of MEM_TREFI : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRCD : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRP : constant is 1;
    attribute mti_svvh_generic_type of MEM_TWR : constant is 1;
    attribute mti_svvh_generic_type of MEM_TWTR : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRTP : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRAS : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRC : constant is 1;
    attribute mti_svvh_generic_type of CFG_TCCD : constant is 1;
    attribute mti_svvh_generic_type of MEM_AUTO_PD_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_RD_TO_WR_TURNAROUND_OCT : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_WR_TO_RD_TURNAROUND_OCT : constant is 1;
    attribute mti_svvh_generic_type of CTL_RD_TO_PCH_EXTRA_CLK : constant is 1;
    attribute mti_svvh_generic_type of CTL_RD_TO_RD_DIFF_CHIP_EXTRA_CLK : constant is 1;
    attribute mti_svvh_generic_type of CTL_WR_TO_WR_DIFF_CHIP_EXTRA_CLK : constant is 1;
    attribute mti_svvh_generic_type of AFI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATE_RATIO : constant is 1;
    attribute mti_svvh_generic_type of AFI_WLAT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RLAT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RRANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_WRANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of USE_SHADOW_REGS : constant is 1;
    attribute mti_svvh_generic_type of CFG_SELF_RFSH_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PDN_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_POWER_SAVING_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_CLK_ENTRY_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of MEM_TMRD_CK : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_AUTO_CORRECTION_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CTL_ECC_MULTIPLES_16_24_40_72 : constant is 1;
    attribute mti_svvh_generic_type of CTL_ENABLE_BURST_INTERRUPT_INT : constant is 1;
    attribute mti_svvh_generic_type of CTL_ENABLE_BURST_TERMINATE_INT : constant is 1;
    attribute mti_svvh_generic_type of CTL_ENABLE_WDATA_PATH_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of CFG_GEN_SBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_GEN_DBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_MASK_SBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_MASK_DBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_MASK_CORRDROP_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_CLR_INTR : constant is 1;
    attribute mti_svvh_generic_type of CTL_USR_REFRESH : constant is 1;
    attribute mti_svvh_generic_type of CTL_REGDIMM_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CFG_WRITE_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_READ_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_WRITE_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_READ_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CKE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_NO_DM : constant is 1;
    attribute mti_svvh_generic_type of CSR_BE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_ERRCMD_FIFO_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_DECODER_REG : constant is 1;
    attribute mti_svvh_generic_type of CTL_CSR_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CSR_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CSR_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ENABLE_BURST_MERGE : constant is 1;
end alt_mem_if_nextgen_ddr2_controller_core;
