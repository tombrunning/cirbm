library verilog;
use verilog.vl_types.all;
entity sequencer_phy_mgr is
    generic(
        AVL_DATA_WIDTH  : integer := 32;
        AVL_ADDR_WIDTH  : integer := 13;
        MAX_LATENCY_COUNT_WIDTH: integer := 5;
        MEM_IF_READ_DQS_WIDTH: integer := 1;
        MEM_IF_WRITE_DQS_WIDTH: integer := 1;
        AFI_DQ_WIDTH    : integer := 64;
        AFI_DEBUG_INFO_WIDTH: integer := 32;
        AFI_MAX_WRITE_LATENCY_COUNT_WIDTH: integer := 5;
        AFI_MAX_READ_LATENCY_COUNT_WIDTH: integer := 5;
        CALIB_VFIFO_OFFSET: integer := 10;
        CALIB_LFIFO_OFFSET: integer := 3;
        CALIB_REG_WIDTH : integer := 8;
        READ_VALID_FIFO_SIZE: integer := 16;
        MEM_T_WL        : integer := 1;
        MEM_T_RL        : integer := 2;
        CTL_REGDIMM_ENABLED: integer := 0;
        NUM_WRITE_FR_CYCLE_SHIFTS: integer := 0;
        DEVICE_FAMILY   : string  := "";
        VFIFO_CONTROL_WIDTH_PER_DQS: integer := 1
    );
    port(
        avl_clk         : in     vl_logic;
        avl_reset_n     : in     vl_logic;
        avl_address     : in     vl_logic_vector;
        avl_write       : in     vl_logic;
        avl_writedata   : in     vl_logic_vector;
        avl_read        : in     vl_logic;
        avl_readdata    : out    vl_logic_vector;
        avl_waitrequest : out    vl_logic;
        phy_clk         : in     vl_logic;
        phy_reset_n     : in     vl_logic;
        phy_read_latency_counter: out    vl_logic_vector;
        phy_read_increment_vfifo_fr: out    vl_logic_vector;
        phy_read_increment_vfifo_hr: out    vl_logic_vector;
        phy_read_increment_vfifo_qr: out    vl_logic_vector;
        phy_reset_mem_stable: out    vl_logic;
        phy_afi_wlat    : out    vl_logic_vector;
        phy_afi_rlat    : out    vl_logic_vector;
        phy_mux_sel     : out    vl_logic;
        phy_cal_success : out    vl_logic;
        phy_cal_fail    : out    vl_logic;
        phy_cal_debug_info: out    vl_logic_vector;
        phy_read_fifo_reset: out    vl_logic_vector;
        phy_vfifo_rd_en_override: out    vl_logic_vector;
        phy_read_fifo_q : in     vl_logic_vector;
        phy_write_fr_cycle_shifts: out    vl_logic_vector;
        calib_skip_steps: in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AVL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AVL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DEBUG_INFO_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_MAX_WRITE_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_MAX_READ_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CALIB_VFIFO_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of CALIB_LFIFO_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of CALIB_REG_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of MEM_T_WL : constant is 1;
    attribute mti_svvh_generic_type of MEM_T_RL : constant is 1;
    attribute mti_svvh_generic_type of CTL_REGDIMM_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of NUM_WRITE_FR_CYCLE_SHIFTS : constant is 1;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of VFIFO_CONTROL_WIDTH_PER_DQS : constant is 1;
end sequencer_phy_mgr;
