library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_s0 is
    port(
        avl_clk         : in     vl_logic;
        avl_reset_n     : in     vl_logic;
        phy_clk         : in     vl_logic;
        phy_reset_n     : in     vl_logic;
        phy_read_latency_counter: out    vl_logic_vector(3 downto 0);
        phy_afi_wlat    : out    vl_logic_vector(5 downto 0);
        phy_afi_rlat    : out    vl_logic_vector(5 downto 0);
        phy_read_increment_vfifo_fr: out    vl_logic_vector(7 downto 0);
        phy_read_increment_vfifo_hr: out    vl_logic_vector(7 downto 0);
        phy_read_increment_vfifo_qr: out    vl_logic_vector(7 downto 0);
        phy_reset_mem_stable: out    vl_logic;
        phy_cal_success : out    vl_logic;
        phy_cal_fail    : out    vl_logic;
        phy_cal_debug_info: out    vl_logic_vector(31 downto 0);
        phy_read_fifo_reset: out    vl_logic_vector(7 downto 0);
        phy_vfifo_rd_en_override: out    vl_logic_vector(7 downto 0);
        phy_read_fifo_q : in     vl_logic_vector(255 downto 0);
        phy_write_fr_cycle_shifts: out    vl_logic_vector(15 downto 0);
        phy_mux_sel     : out    vl_logic;
        calib_skip_steps: in     vl_logic_vector(7 downto 0);
        afi_clk         : in     vl_logic;
        afi_reset_n     : in     vl_logic;
        afi_addr        : out    vl_logic_vector(27 downto 0);
        afi_ba          : out    vl_logic_vector(5 downto 0);
        afi_cs_n        : out    vl_logic_vector(1 downto 0);
        afi_cke         : out    vl_logic_vector(1 downto 0);
        afi_odt         : out    vl_logic_vector(1 downto 0);
        afi_ras_n       : out    vl_logic_vector(1 downto 0);
        afi_cas_n       : out    vl_logic_vector(1 downto 0);
        afi_we_n        : out    vl_logic_vector(1 downto 0);
        afi_dqs_burst   : out    vl_logic_vector(15 downto 0);
        afi_wdata       : out    vl_logic_vector(255 downto 0);
        afi_wdata_valid : out    vl_logic_vector(15 downto 0);
        afi_dm          : out    vl_logic_vector(31 downto 0);
        afi_rdata_en    : out    vl_logic_vector(1 downto 0);
        afi_rdata_en_full: out    vl_logic_vector(1 downto 0);
        afi_rdata       : in     vl_logic_vector(255 downto 0);
        afi_rdata_valid : in     vl_logic_vector(1 downto 0);
        scc_data        : out    vl_logic;
        scc_dqs_ena     : out    vl_logic_vector(7 downto 0);
        scc_dqs_io_ena  : out    vl_logic_vector(7 downto 0);
        scc_dq_ena      : out    vl_logic_vector(63 downto 0);
        scc_dm_ena      : out    vl_logic_vector(7 downto 0);
        capture_strobe_tracking: in     vl_logic_vector(7 downto 0);
        scc_upd         : out    vl_logic_vector(0 downto 0);
        afi_init_req    : in     vl_logic;
        afi_cal_req     : in     vl_logic;
        scc_clk         : in     vl_logic;
        reset_n_scc_clk : in     vl_logic
    );
end DE4_QSYS_mem_if_ddr2_emif_s0;
