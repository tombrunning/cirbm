library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_timing_param is
    generic(
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_CTL_ARBITER_TYPE: string  := "ROWCOL";
        CFG_PORT_WIDTH_TYPE: integer := 3;
        CFG_PORT_WIDTH_BURST_LENGTH: integer := 5;
        CFG_PORT_WIDTH_CAS_WR_LAT: integer := 4;
        CFG_PORT_WIDTH_ADD_LAT: integer := 3;
        CFG_PORT_WIDTH_TCL: integer := 4;
        CFG_PORT_WIDTH_TRRD: integer := 4;
        CFG_PORT_WIDTH_TFAW: integer := 6;
        CFG_PORT_WIDTH_TRFC: integer := 8;
        CFG_PORT_WIDTH_TREFI: integer := 13;
        CFG_PORT_WIDTH_TRCD: integer := 4;
        CFG_PORT_WIDTH_TRP: integer := 4;
        CFG_PORT_WIDTH_TWR: integer := 4;
        CFG_PORT_WIDTH_TWTR: integer := 4;
        CFG_PORT_WIDTH_TRTP: integer := 4;
        CFG_PORT_WIDTH_TRAS: integer := 5;
        CFG_PORT_WIDTH_TRC: integer := 6;
        CFG_PORT_WIDTH_TCCD: integer := 3;
        CFG_PORT_WIDTH_TMRD: integer := 3;
        CFG_PORT_WIDTH_SELF_RFSH_EXIT_CYCLES: integer := 10;
        CFG_PORT_WIDTH_PDN_EXIT_CYCLES: integer := 4;
        CFG_PORT_WIDTH_AUTO_PD_CYCLES: integer := 16;
        CFG_PORT_WIDTH_POWER_SAVING_EXIT_CYCLES: integer := 4;
        CFG_PORT_WIDTH_MEM_CLK_ENTRY_CYCLES: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_RDWR: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_PCH: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_BC: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_PCH: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_AP_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_BC: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_PCH: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_AP_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_ALL_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT_DIFF_BANK: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_FOUR_ACT_TO_ACT: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_ZQ_CAL: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_PERIOD: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_PERIOD: integer := 4;
        T_PARAM_ACT_TO_RDWR_WIDTH: integer := 6;
        T_PARAM_ACT_TO_PCH_WIDTH: integer := 6;
        T_PARAM_ACT_TO_ACT_WIDTH: integer := 6;
        T_PARAM_RD_TO_RD_WIDTH: integer := 6;
        T_PARAM_RD_TO_RD_DIFF_CHIP_WIDTH: integer := 6;
        T_PARAM_RD_TO_WR_WIDTH: integer := 6;
        T_PARAM_RD_TO_WR_BC_WIDTH: integer := 6;
        T_PARAM_RD_TO_WR_DIFF_CHIP_WIDTH: integer := 6;
        T_PARAM_RD_TO_PCH_WIDTH: integer := 6;
        T_PARAM_RD_AP_TO_VALID_WIDTH: integer := 6;
        T_PARAM_WR_TO_WR_WIDTH: integer := 6;
        T_PARAM_WR_TO_WR_DIFF_CHIP_WIDTH: integer := 6;
        T_PARAM_WR_TO_RD_WIDTH: integer := 6;
        T_PARAM_WR_TO_RD_BC_WIDTH: integer := 6;
        T_PARAM_WR_TO_RD_DIFF_CHIP_WIDTH: integer := 6;
        T_PARAM_WR_TO_PCH_WIDTH: integer := 6;
        T_PARAM_WR_AP_TO_VALID_WIDTH: integer := 6;
        T_PARAM_PCH_TO_VALID_WIDTH: integer := 6;
        T_PARAM_PCH_ALL_TO_VALID_WIDTH: integer := 6;
        T_PARAM_ACT_TO_ACT_DIFF_BANK_WIDTH: integer := 6;
        T_PARAM_FOUR_ACT_TO_ACT_WIDTH: integer := 6;
        T_PARAM_ARF_TO_VALID_WIDTH: integer := 8;
        T_PARAM_PDN_TO_VALID_WIDTH: integer := 6;
        T_PARAM_SRF_TO_VALID_WIDTH: integer := 10;
        T_PARAM_SRF_TO_ZQ_CAL_WIDTH: integer := 10;
        T_PARAM_ARF_PERIOD_WIDTH: integer := 13;
        T_PARAM_PDN_PERIOD_WIDTH: integer := 16;
        T_PARAM_POWER_SAVING_EXIT_WIDTH: integer := 6;
        T_PARAM_MEM_CLK_ENTRY_CYCLES_WIDTH: integer := 4
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        cfg_burst_length: in     vl_logic_vector;
        cfg_type        : in     vl_logic_vector;
        cfg_cas_wr_lat  : in     vl_logic_vector;
        cfg_add_lat     : in     vl_logic_vector;
        cfg_tcl         : in     vl_logic_vector;
        cfg_trrd        : in     vl_logic_vector;
        cfg_tfaw        : in     vl_logic_vector;
        cfg_trfc        : in     vl_logic_vector;
        cfg_trefi       : in     vl_logic_vector;
        cfg_trcd        : in     vl_logic_vector;
        cfg_trp         : in     vl_logic_vector;
        cfg_twr         : in     vl_logic_vector;
        cfg_twtr        : in     vl_logic_vector;
        cfg_trtp        : in     vl_logic_vector;
        cfg_tras        : in     vl_logic_vector;
        cfg_trc         : in     vl_logic_vector;
        cfg_tccd        : in     vl_logic_vector;
        cfg_tmrd        : in     vl_logic_vector;
        cfg_self_rfsh_exit_cycles: in     vl_logic_vector;
        cfg_pdn_exit_cycles: in     vl_logic_vector;
        cfg_auto_pd_cycles: in     vl_logic_vector;
        cfg_power_saving_exit_cycles: in     vl_logic_vector;
        cfg_mem_clk_entry_cycles: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_rdwr: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_pch: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_act: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_rd: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_rd_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_wr: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_wr_bc: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_wr_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_pch: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_ap_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_wr: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_wr_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_rd: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_rd_bc: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_rd_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_pch: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_ap_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_pch_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_pch_all_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_act_diff_bank: in     vl_logic_vector;
        cfg_extra_ctl_clk_four_act_to_act: in     vl_logic_vector;
        cfg_extra_ctl_clk_arf_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_pdn_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_srf_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_srf_to_zq_cal: in     vl_logic_vector;
        cfg_extra_ctl_clk_arf_period: in     vl_logic_vector;
        cfg_extra_ctl_clk_pdn_period: in     vl_logic_vector;
        t_param_act_to_rdwr: out    vl_logic_vector;
        t_param_act_to_pch: out    vl_logic_vector;
        t_param_act_to_act: out    vl_logic_vector;
        t_param_rd_to_rd: out    vl_logic_vector;
        t_param_rd_to_rd_diff_chip: out    vl_logic_vector;
        t_param_rd_to_wr: out    vl_logic_vector;
        t_param_rd_to_wr_bc: out    vl_logic_vector;
        t_param_rd_to_wr_diff_chip: out    vl_logic_vector;
        t_param_rd_to_pch: out    vl_logic_vector;
        t_param_rd_ap_to_valid: out    vl_logic_vector;
        t_param_wr_to_wr: out    vl_logic_vector;
        t_param_wr_to_wr_diff_chip: out    vl_logic_vector;
        t_param_wr_to_rd: out    vl_logic_vector;
        t_param_wr_to_rd_bc: out    vl_logic_vector;
        t_param_wr_to_rd_diff_chip: out    vl_logic_vector;
        t_param_wr_to_pch: out    vl_logic_vector;
        t_param_wr_ap_to_valid: out    vl_logic_vector;
        t_param_pch_to_valid: out    vl_logic_vector;
        t_param_pch_all_to_valid: out    vl_logic_vector;
        t_param_act_to_act_diff_bank: out    vl_logic_vector;
        t_param_four_act_to_act: out    vl_logic_vector;
        t_param_arf_to_valid: out    vl_logic_vector;
        t_param_pdn_to_valid: out    vl_logic_vector;
        t_param_srf_to_valid: out    vl_logic_vector;
        t_param_srf_to_zq_cal: out    vl_logic_vector;
        t_param_arf_period: out    vl_logic_vector;
        t_param_pdn_period: out    vl_logic_vector;
        t_param_power_saving_exit: out    vl_logic_vector;
        t_param_mem_clk_entry_cycles: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_CTL_ARBITER_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_BURST_LENGTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_CAS_WR_LAT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ADD_LAT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TCL : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRRD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TFAW : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRFC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TREFI : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRCD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TWR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TWTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRTP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRAS : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TCCD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TMRD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_SELF_RFSH_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_PDN_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_AUTO_PD_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_POWER_SAVING_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MEM_CLK_ENTRY_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_RDWR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_PCH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_BC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_PCH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_AP_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_BC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_PCH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_AP_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_ALL_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT_DIFF_BANK : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_FOUR_ACT_TO_ACT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_ZQ_CAL : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_RDWR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_PCH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_ACT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_RD_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_RD_DIFF_CHIP_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_WR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_WR_BC_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_WR_DIFF_CHIP_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_PCH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_AP_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_WR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_WR_DIFF_CHIP_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_RD_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_RD_BC_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_RD_DIFF_CHIP_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_PCH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_AP_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_PCH_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_PCH_ALL_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_ACT_DIFF_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_FOUR_ACT_TO_ACT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ARF_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_PDN_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_SRF_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_SRF_TO_ZQ_CAL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ARF_PERIOD_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_PDN_PERIOD_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_POWER_SAVING_EXIT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_MEM_CLK_ENTRY_CYCLES_WIDTH : constant is 1;
end alt_mem_ddrx_timing_param;
