library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_rdwr_data_tmg is
    generic(
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_MEM_IF_CHIP : integer := 1;
        CFG_MEM_IF_DQ_WIDTH: integer := 8;
        CFG_MEM_IF_DQS_WIDTH: integer := 1;
        CFG_MEM_IF_DM_WIDTH: integer := 1;
        CFG_WLAT_BUS_WIDTH: integer := 6;
        CFG_DRAM_WLAT_GROUP: integer := 1;
        CFG_DATA_ID_WIDTH: integer := 10;
        CFG_WDATA_REG   : integer := 0;
        CFG_ECC_ENC_REG : integer := 0;
        CFG_AFI_INTF_PHASE_NUM: integer := 2;
        CFG_PORT_WIDTH_ENABLE_ECC: integer := 1;
        CFG_PORT_WIDTH_OUTPUT_REGD: integer := 1;
        CFG_CTL_ARBITER_TYPE: string  := "ROWCOL";
        CFG_USE_SHADOW_REGS: integer := 0
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        cfg_enable_ecc  : in     vl_logic_vector;
        cfg_output_regd : in     vl_logic_vector;
        cfg_output_regd_for_afi_output: out    vl_logic_vector;
        bg_do_read      : in     vl_logic_vector;
        bg_do_write     : in     vl_logic_vector;
        bg_doing_read   : in     vl_logic;
        bg_doing_write  : in     vl_logic;
        bg_rdwr_data_valid: in     vl_logic;
        dataid          : in     vl_logic_vector;
        bg_do_rmw_correct: in     vl_logic_vector;
        bg_do_rmw_partial: in     vl_logic_vector;
        bg_to_chip      : in     vl_logic_vector;
        ecc_wdata       : in     vl_logic_vector;
        ecc_dm          : in     vl_logic_vector;
        afi_wlat        : in     vl_logic_vector;
        afi_doing_read  : out    vl_logic_vector;
        afi_doing_read_full: out    vl_logic_vector;
        ecc_wdata_fifo_read: out    vl_logic_vector;
        ecc_wdata_fifo_dataid: out    vl_logic_vector;
        ecc_wdata_fifo_dataid_vector: out    vl_logic_vector;
        ecc_wdata_fifo_rmw_correct: out    vl_logic_vector;
        ecc_wdata_fifo_rmw_partial: out    vl_logic_vector;
        ecc_wdata_fifo_read_first: out    vl_logic;
        ecc_wdata_fifo_dataid_first: out    vl_logic_vector;
        ecc_wdata_fifo_dataid_vector_first: out    vl_logic_vector;
        ecc_wdata_fifo_rmw_correct_first: out    vl_logic;
        ecc_wdata_fifo_rmw_partial_first: out    vl_logic;
        ecc_wdata_fifo_first_vector: out    vl_logic_vector;
        ecc_wdata_fifo_read_last: out    vl_logic;
        ecc_wdata_fifo_dataid_last: out    vl_logic_vector;
        ecc_wdata_fifo_dataid_vector_last: out    vl_logic_vector;
        ecc_wdata_fifo_rmw_correct_last: out    vl_logic;
        ecc_wdata_fifo_rmw_partial_last: out    vl_logic;
        afi_rrank       : out    vl_logic_vector;
        afi_wrank       : out    vl_logic_vector;
        afi_dqs_burst   : out    vl_logic_vector;
        afi_wdata_valid : out    vl_logic_vector;
        afi_wdata       : out    vl_logic_vector;
        afi_dm          : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_WLAT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DRAM_WLAT_GROUP : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_WDATA_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_ENC_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_AFI_INTF_PHASE_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_ECC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_OUTPUT_REGD : constant is 1;
    attribute mti_svvh_generic_type of CFG_CTL_ARBITER_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_USE_SHADOW_REGS : constant is 1;
end alt_mem_ddrx_rdwr_data_tmg;
