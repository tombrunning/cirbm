library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_wdata_path is
    generic(
        CFG_LOCAL_DATA_WIDTH: integer := 16;
        CFG_MEM_IF_DQ_WIDTH: integer := 8;
        CFG_MEM_IF_DQS_WIDTH: integer := 1;
        CFG_INT_SIZE_WIDTH: integer := 5;
        CFG_DATA_ID_WIDTH: integer := 4;
        CFG_DRAM_WLAT_GROUP: integer := 1;
        CFG_LOCAL_WLAT_GROUP: integer := 1;
        CFG_TBP_NUM     : integer := 8;
        CFG_BUFFER_ADDR_WIDTH: integer := 10;
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_ECC_MULTIPLES: integer := 1;
        CFG_WDATA_REG   : integer := 0;
        CFG_PARTIAL_BE_PER_WORD_ENABLE: integer := 1;
        CFG_ECC_CODE_WIDTH: integer := 8;
        CFG_PORT_WIDTH_BURST_LENGTH: integer := 5;
        CFG_PORT_WIDTH_ENABLE_ECC: integer := 1;
        CFG_PORT_WIDTH_ENABLE_AUTO_CORR: integer := 1;
        CFG_PORT_WIDTH_ENABLE_NO_DM: integer := 1;
        CFG_PORT_WIDTH_ENABLE_ECC_CODE_OVERWRITES: integer := 1;
        CFG_PORT_WIDTH_INTERFACE_WIDTH: integer := 8
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        cfg_burst_length: in     vl_logic_vector;
        cfg_enable_ecc  : in     vl_logic_vector;
        cfg_enable_auto_corr: in     vl_logic_vector;
        cfg_enable_no_dm: in     vl_logic_vector;
        cfg_enable_ecc_code_overwrites: in     vl_logic_vector;
        cfg_interface_width: in     vl_logic_vector;
        wdatap_free_id_valid: out    vl_logic;
        wdatap_free_id_dataid: out    vl_logic_vector;
        proc_busy       : in     vl_logic;
        proc_load       : in     vl_logic;
        proc_load_dataid: in     vl_logic;
        proc_write      : in     vl_logic;
        tbp_load_index  : in     vl_logic_vector;
        proc_size       : in     vl_logic_vector;
        wr_data_mem_full: out    vl_logic;
        write_data_en   : in     vl_logic;
        write_data      : in     vl_logic_vector;
        byte_en         : in     vl_logic_vector;
        data_complete   : out    vl_logic_vector;
        data_rmw_complete: out    vl_logic;
        data_rmw_fetch  : in     vl_logic;
        data_partial_be : out    vl_logic;
        doing_write     : in     vl_logic_vector;
        dataid          : in     vl_logic_vector;
        dataid_vector   : in     vl_logic_vector;
        rdwr_data_valid : in     vl_logic_vector;
        rmw_correct     : in     vl_logic_vector;
        rmw_partial     : in     vl_logic_vector;
        doing_write_first: in     vl_logic;
        dataid_first    : in     vl_logic_vector;
        dataid_vector_first: in     vl_logic_vector;
        rdwr_data_valid_first: in     vl_logic;
        rmw_correct_first: in     vl_logic;
        rmw_partial_first: in     vl_logic;
        doing_write_first_vector: in     vl_logic_vector;
        rdwr_data_valid_first_vector: in     vl_logic_vector;
        doing_write_last: in     vl_logic;
        dataid_last     : in     vl_logic_vector;
        dataid_vector_last: in     vl_logic_vector;
        rdwr_data_valid_last: in     vl_logic;
        rmw_correct_last: in     vl_logic;
        rmw_partial_last: in     vl_logic;
        wdatap_data     : out    vl_logic_vector;
        wdatap_rmw_partial_data: out    vl_logic_vector;
        wdatap_rmw_correct_data: out    vl_logic_vector;
        wdatap_rmw_partial: out    vl_logic;
        wdatap_rmw_correct: out    vl_logic;
        wdatap_dm       : out    vl_logic_vector;
        wdatap_ecc_code : out    vl_logic_vector;
        wdatap_ecc_code_overwrite: out    vl_logic_vector;
        rmwfifo_data_valid: in     vl_logic;
        rmwfifo_data    : in     vl_logic_vector;
        rmwfifo_ecc_dbe : in     vl_logic_vector;
        rmwfifo_ecc_code: in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_INT_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DRAM_WLAT_GROUP : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_WLAT_GROUP : constant is 1;
    attribute mti_svvh_generic_type of CFG_TBP_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_BUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_MULTIPLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_WDATA_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_PARTIAL_BE_PER_WORD_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_CODE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_BURST_LENGTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_ECC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_AUTO_CORR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_NO_DM : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_ECC_CODE_OVERWRITES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_INTERFACE_WIDTH : constant is 1;
end alt_mem_ddrx_wdata_path;
