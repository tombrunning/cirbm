library verilog;
use verilog.vl_types.all;
entity rw_manager_ddr2 is
    generic(
        AVL_DATA_WIDTH  : integer := 32;
        AVL_ADDR_WIDTH  : integer := 16;
        MEM_ADDRESS_WIDTH: integer := 19;
        MEM_CONTROL_WIDTH: integer := 4;
        MEM_DQ_WIDTH    : integer := 36;
        MEM_DM_WIDTH    : integer := 4;
        MEM_NUMBER_OF_RANKS: integer := 1;
        MEM_CLK_EN_WIDTH: integer := 1;
        MEM_BANK_WIDTH  : integer := 2;
        MEM_ODT_WIDTH   : integer := 1;
        MEM_CHIP_SELECT_WIDTH: integer := 1;
        MEM_READ_DQS_WIDTH: integer := 4;
        MEM_WRITE_DQS_WIDTH: integer := 4;
        AFI_RATIO       : integer := 2;
        RATE            : string  := "Half";
        HCX_COMPAT_MODE : integer := 0;
        DEVICE_FAMILY   : string  := "STRATIXIV";
        AC_ROM_INIT_FILE_NAME: string  := "AC_ROM.hex";
        INST_ROM_INIT_FILE_NAME: string  := "inst_ROM.hex";
        DEBUG_WRITE_TO_READ_RATIO_2_EXPONENT: integer := 0;
        DEBUG_WRITE_TO_READ_RATIO: integer := 0;
        MAX_DI_BUFFER_WORDS_LOG_2: integer := 0;
        AC_BUS_WIDTH    : integer := 30
    );
    port(
        avl_clk         : in     vl_logic;
        avl_reset_n     : in     vl_logic;
        avl_address     : in     vl_logic_vector;
        avl_write       : in     vl_logic;
        avl_writedata   : in     vl_logic_vector;
        avl_read        : in     vl_logic;
        avl_readdata    : out    vl_logic_vector;
        avl_waitrequest : out    vl_logic;
        afi_clk         : in     vl_logic;
        afi_reset_n     : in     vl_logic;
        afi_addr        : out    vl_logic_vector;
        afi_ba          : out    vl_logic_vector;
        afi_cs_n        : out    vl_logic_vector;
        afi_cke         : out    vl_logic_vector;
        afi_odt         : out    vl_logic_vector;
        afi_ras_n       : out    vl_logic_vector;
        afi_cas_n       : out    vl_logic_vector;
        afi_we_n        : out    vl_logic_vector;
        afi_dqs_burst   : out    vl_logic_vector;
        afi_wdata       : out    vl_logic_vector;
        afi_wdata_valid : out    vl_logic_vector;
        afi_dm          : out    vl_logic_vector;
        afi_rdata_en    : out    vl_logic_vector;
        afi_rdata_en_full: out    vl_logic_vector;
        afi_rdata       : in     vl_logic_vector;
        afi_rdata_valid : in     vl_logic_vector;
        csr_clk         : in     vl_logic;
        csr_ena         : in     vl_logic;
        csr_dout_phy    : in     vl_logic;
        csr_dout        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AVL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AVL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_NUMBER_OF_RANKS : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CHIP_SELECT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATIO : constant is 1;
    attribute mti_svvh_generic_type of RATE : constant is 1;
    attribute mti_svvh_generic_type of HCX_COMPAT_MODE : constant is 1;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of AC_ROM_INIT_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of INST_ROM_INIT_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_WRITE_TO_READ_RATIO_2_EXPONENT : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_WRITE_TO_READ_RATIO : constant is 1;
    attribute mti_svvh_generic_type of MAX_DI_BUFFER_WORDS_LOG_2 : constant is 1;
    attribute mti_svvh_generic_type of AC_BUS_WIDTH : constant is 1;
end rw_manager_ddr2;
