library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_p0_read_datapath is
    generic(
        DEVICE_FAMILY   : string  := "";
        MEM_ADDRESS_WIDTH: string  := "";
        MEM_DM_WIDTH    : string  := "";
        MEM_CONTROL_WIDTH: string  := "";
        MEM_DQ_WIDTH    : string  := "";
        MEM_READ_DQS_WIDTH: string  := "";
        MEM_WRITE_DQS_WIDTH: string  := "";
        AFI_ADDRESS_WIDTH: string  := "";
        AFI_DATA_MASK_WIDTH: string  := "";
        AFI_CONTROL_WIDTH: string  := "";
        AFI_DATA_WIDTH  : string  := "";
        AFI_DQS_WIDTH   : string  := "";
        AFI_RATE_RATIO  : string  := "";
        MAX_LATENCY_COUNT_WIDTH: string  := "";
        MAX_READ_LATENCY: string  := "";
        READ_FIFO_READ_MEM_DEPTH: string  := "";
        READ_FIFO_READ_ADDR_WIDTH: string  := "";
        READ_FIFO_WRITE_MEM_DEPTH: string  := "";
        READ_FIFO_WRITE_ADDR_WIDTH: string  := "";
        READ_VALID_FIFO_SIZE: string  := "";
        READ_VALID_FIFO_READ_MEM_DEPTH: string  := "";
        READ_VALID_FIFO_READ_ADDR_WIDTH: string  := "";
        READ_VALID_FIFO_WRITE_MEM_DEPTH: string  := "";
        READ_VALID_FIFO_WRITE_ADDR_WIDTH: string  := "";
        READ_VALID_FIFO_PER_DQS_WIDTH: string  := "";
        NUM_SUBGROUP_PER_READ_DQS: string  := "";
        MEM_T_RL        : string  := "";
        QVLD_EXTRA_FLOP_STAGES: string  := "";
        QVLD_WR_ADDRESS_OFFSET: string  := "";
        REGISTER_C2P    : string  := "";
        VFIFO_C2P_PIPELINE_DEPTH: integer := 1;
        CALIB_REG_WIDTH : string  := "";
        FAST_SIM_MODEL  : string  := "";
        EXTRA_VFIFO_SHIFT: integer := 0
    );
    port(
        reset_n_afi_clk : in     vl_logic;
        seq_read_fifo_reset: in     vl_logic_vector;
        reset_n_resync_clk: in     vl_logic;
        pll_dqs_ena_clk : in     vl_logic;
        read_capture_clk: in     vl_logic_vector;
        ddio_phy_dq     : in     vl_logic_vector;
        pll_afi_clk     : in     vl_logic;
        seq_read_latency_counter: in     vl_logic_vector;
        seq_read_increment_vfifo_fr: in     vl_logic_vector;
        seq_read_increment_vfifo_hr: in     vl_logic_vector;
        seq_read_increment_vfifo_qr: in     vl_logic_vector;
        afi_rdata_en    : in     vl_logic_vector;
        afi_rdata_en_full: in     vl_logic_vector;
        afi_rdata       : out    vl_logic_vector;
        phy_mux_read_fifo_q: out    vl_logic_vector;
        force_oct_off   : out    vl_logic_vector;
        dqs_enable_ctrl : out    vl_logic_vector;
        afi_rdata_valid : out    vl_logic_vector;
        seq_calib_init  : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DATA_MASK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATE_RATIO : constant is 1;
    attribute mti_svvh_generic_type of MAX_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_READ_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of READ_FIFO_READ_MEM_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of READ_FIFO_READ_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of READ_FIFO_WRITE_MEM_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of READ_FIFO_WRITE_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_READ_MEM_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_READ_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_WRITE_MEM_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_WRITE_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_PER_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_SUBGROUP_PER_READ_DQS : constant is 1;
    attribute mti_svvh_generic_type of MEM_T_RL : constant is 1;
    attribute mti_svvh_generic_type of QVLD_EXTRA_FLOP_STAGES : constant is 1;
    attribute mti_svvh_generic_type of QVLD_WR_ADDRESS_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of REGISTER_C2P : constant is 1;
    attribute mti_svvh_generic_type of VFIFO_C2P_PIPELINE_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of CALIB_REG_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of FAST_SIM_MODEL : constant is 1;
    attribute mti_svvh_generic_type of EXTRA_VFIFO_SHIFT : constant is 1;
end DE4_QSYS_mem_if_ddr2_emif_p0_read_datapath;
