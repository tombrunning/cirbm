library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_controller is
    generic(
        CFG_LOCAL_SIZE_WIDTH: integer := 3;
        CFG_LOCAL_ADDR_WIDTH: integer := 32;
        CFG_LOCAL_DATA_WIDTH: integer := 80;
        CFG_LOCAL_ID_WIDTH: integer := 8;
        CFG_LOCAL_IF_TYPE: string  := "AVALON";
        CFG_MEM_IF_CHIP : integer := 2;
        CFG_MEM_IF_CS_WIDTH: integer := 1;
        CFG_MEM_IF_BA_WIDTH: integer := 3;
        CFG_MEM_IF_ROW_WIDTH: integer := 15;
        CFG_MEM_IF_COL_WIDTH: integer := 12;
        CFG_MEM_IF_ADDR_WIDTH: integer := 15;
        CFG_MEM_IF_CKE_WIDTH: integer := 2;
        CFG_MEM_IF_ODT_WIDTH: integer := 2;
        CFG_MEM_IF_CLK_PAIR_COUNT: integer := 2;
        CFG_MEM_IF_DQ_WIDTH: integer := 40;
        CFG_MEM_IF_DQS_WIDTH: integer := 5;
        CFG_MEM_IF_DM_WIDTH: integer := 5;
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_ODT_ENABLED : integer := 1;
        \CFG_OUTPUT_REGD\: integer := 0;
        CFG_CTL_TBP_NUM : integer := 4;
        CFG_LPDDR2_ENABLED: integer := 0;
        CFG_DATA_REORDERING_TYPE: string  := "INTER_BANK";
        CFG_ECC_MULTIPLES_16_24_40_72: integer := 1;
        CFG_WRBUFFER_ADDR_WIDTH: integer := 6;
        CFG_RDBUFFER_ADDR_WIDTH: integer := 10;
        CFG_MAX_PENDING_RD_CMD: integer := 16;
        CFG_MAX_PENDING_WR_CMD: integer := 8;
        CFG_PORT_WIDTH_TYPE: integer := 3;
        CFG_PORT_WIDTH_INTERFACE_WIDTH: integer := 8;
        CFG_PORT_WIDTH_BURST_LENGTH: integer := 5;
        CFG_PORT_WIDTH_DEVICE_WIDTH: integer := 4;
        CFG_PORT_WIDTH_OUTPUT_REGD: integer := 2;
        CFG_PORT_WIDTH_ADDR_ORDER: integer := 2;
        CFG_PORT_WIDTH_COL_ADDR_WIDTH: integer := 5;
        CFG_PORT_WIDTH_ROW_ADDR_WIDTH: integer := 5;
        CFG_PORT_WIDTH_BANK_ADDR_WIDTH: integer := 3;
        CFG_PORT_WIDTH_CS_ADDR_WIDTH: integer := 3;
        CFG_PORT_WIDTH_CAS_WR_LAT: integer := 4;
        CFG_PORT_WIDTH_ADD_LAT: integer := 3;
        CFG_PORT_WIDTH_TCL: integer := 4;
        CFG_PORT_WIDTH_TRRD: integer := 4;
        CFG_PORT_WIDTH_TFAW: integer := 6;
        CFG_PORT_WIDTH_TRFC: integer := 8;
        CFG_PORT_WIDTH_TREFI: integer := 13;
        CFG_PORT_WIDTH_TRCD: integer := 4;
        CFG_PORT_WIDTH_TRP: integer := 4;
        CFG_PORT_WIDTH_TWR: integer := 4;
        CFG_PORT_WIDTH_TWTR: integer := 4;
        CFG_PORT_WIDTH_TRTP: integer := 4;
        CFG_PORT_WIDTH_TRAS: integer := 5;
        CFG_PORT_WIDTH_TRC: integer := 6;
        CFG_PORT_WIDTH_TCCD: integer := 4;
        CFG_PORT_WIDTH_TMRD: integer := 3;
        CFG_PORT_WIDTH_SELF_RFSH_EXIT_CYCLES: integer := 10;
        CFG_PORT_WIDTH_PDN_EXIT_CYCLES: integer := 4;
        CFG_PORT_WIDTH_AUTO_PD_CYCLES: integer := 16;
        CFG_PORT_WIDTH_POWER_SAVING_EXIT_CYCLES: integer := 4;
        CFG_PORT_WIDTH_MEM_CLK_ENTRY_CYCLES: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_RDWR: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_PCH: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_BC: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_PCH: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_AP_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_BC: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_DIFF_CHIP: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_PCH: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_AP_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_ALL_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT_DIFF_BANK: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_FOUR_ACT_TO_ACT: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_VALID: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_ZQ_CAL: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_PERIOD: integer := 4;
        CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_PERIOD: integer := 4;
        CFG_PORT_WIDTH_REORDER_DATA: integer := 1;
        CFG_PORT_WIDTH_STARVE_LIMIT: integer := 6;
        CFG_PORT_WIDTH_USER_RFSH: integer := 1;
        CFG_PORT_WIDTH_SELF_RFSH: integer := 1;
        CFG_PORT_WIDTH_REGDIMM_ENABLE: integer := 1;
        CFG_PORT_WIDTH_ENABLE_BURST_INTERRUPT: integer := 1;
        CFG_PORT_WIDTH_ENABLE_BURST_TERMINATE: integer := 1;
        CFG_ENABLE_CMD_SPLIT: vl_logic := Hi1;
        CFG_ENABLE_WDATA_PATH_LATENCY: integer := 0;
        CFG_PORT_WIDTH_ENABLE_ECC: integer := 1;
        CFG_PORT_WIDTH_ENABLE_AUTO_CORR: integer := 1;
        CFG_PORT_WIDTH_GEN_SBE: integer := 1;
        CFG_PORT_WIDTH_GEN_DBE: integer := 1;
        CFG_PORT_WIDTH_ENABLE_INTR: integer := 1;
        CFG_PORT_WIDTH_MASK_SBE_INTR: integer := 1;
        CFG_PORT_WIDTH_MASK_DBE_INTR: integer := 1;
        CFG_PORT_WIDTH_MASK_CORR_DROPPED_INTR: integer := 1;
        CFG_PORT_WIDTH_CLR_INTR: integer := 1;
        CFG_PORT_WIDTH_ENABLE_ECC_CODE_OVERWRITES: integer := 1;
        CFG_PORT_WIDTH_ENABLE_NO_DM: integer := 1;
        CFG_ECC_DECODER_REG: integer := 1;
        CFG_PORT_WIDTH_WRITE_ODT_CHIP: integer := 4;
        CFG_PORT_WIDTH_READ_ODT_CHIP: integer := 4;
        STS_PORT_WIDTH_SBE_ERROR: integer := 1;
        STS_PORT_WIDTH_DBE_ERROR: integer := 1;
        STS_PORT_WIDTH_CORR_DROP_ERROR: integer := 1;
        STS_PORT_WIDTH_SBE_COUNT: integer := 8;
        STS_PORT_WIDTH_DBE_COUNT: integer := 8;
        STS_PORT_WIDTH_CORR_DROP_COUNT: integer := 8;
        CFG_WLAT_BUS_WIDTH: integer := 4;
        CFG_RRANK_BUS_WIDTH: integer := 1;
        CFG_WRANK_BUS_WIDTH: integer := 1;
        CFG_USE_SHADOW_REGS: integer := 0;
        CFG_RDATA_RETURN_MODE: string  := "PASSTHROUGH";
        CFG_ERRCMD_FIFO_REG: integer := 0;
        CFG_ENABLE_BURST_MERGE: integer := 0
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        itf_cmd_ready   : out    vl_logic;
        itf_cmd_valid   : in     vl_logic;
        itf_cmd         : in     vl_logic;
        itf_cmd_address : in     vl_logic_vector;
        itf_cmd_burstlen: in     vl_logic_vector;
        itf_cmd_id      : in     vl_logic_vector;
        itf_cmd_priority: in     vl_logic;
        itf_cmd_autopercharge: in     vl_logic;
        itf_cmd_multicast: in     vl_logic;
        itf_wr_data_ready: out    vl_logic;
        itf_wr_data_valid: in     vl_logic;
        itf_wr_data     : in     vl_logic_vector;
        itf_wr_data_byte_en: in     vl_logic_vector;
        itf_wr_data_begin: in     vl_logic;
        itf_wr_data_last: in     vl_logic;
        itf_wr_data_id  : in     vl_logic_vector;
        itf_rd_data_ready: in     vl_logic;
        itf_rd_data_valid: out    vl_logic;
        itf_rd_data     : out    vl_logic_vector;
        itf_rd_data_error: out    vl_logic;
        itf_rd_data_begin: out    vl_logic;
        itf_rd_data_last: out    vl_logic;
        itf_rd_data_id  : out    vl_logic_vector;
        itf_rd_data_id_early: out    vl_logic_vector;
        itf_rd_data_id_early_valid: out    vl_logic;
        local_refresh_req: in     vl_logic;
        local_refresh_chip: in     vl_logic_vector;
        local_zqcal_req : in     vl_logic;
        local_zqcal_chip: in     vl_logic_vector;
        local_deep_powerdn_chip: in     vl_logic_vector;
        local_deep_powerdn_req: in     vl_logic;
        local_self_rfsh_req: in     vl_logic;
        local_self_rfsh_chip: in     vl_logic_vector;
        local_refresh_ack: out    vl_logic;
        local_deep_powerdn_ack: out    vl_logic;
        local_power_down_ack: out    vl_logic;
        local_self_rfsh_ack: out    vl_logic;
        local_init_done : out    vl_logic;
        afi_rst_n       : out    vl_logic_vector;
        afi_ba          : out    vl_logic_vector;
        afi_addr        : out    vl_logic_vector;
        afi_cke         : out    vl_logic_vector;
        afi_cs_n        : out    vl_logic_vector;
        afi_ras_n       : out    vl_logic_vector;
        afi_cas_n       : out    vl_logic_vector;
        afi_we_n        : out    vl_logic_vector;
        afi_odt         : out    vl_logic_vector;
        afi_wlat        : in     vl_logic_vector;
        afi_dqs_burst   : out    vl_logic_vector;
        afi_dm          : out    vl_logic_vector;
        afi_wdata       : out    vl_logic_vector;
        afi_wdata_valid : out    vl_logic_vector;
        afi_rdata_en    : out    vl_logic_vector;
        afi_rdata_en_full: out    vl_logic_vector;
        afi_rrank       : out    vl_logic_vector;
        afi_wrank       : out    vl_logic_vector;
        afi_rdata       : in     vl_logic_vector;
        afi_rdata_valid : in     vl_logic_vector;
        ctl_cal_success : in     vl_logic;
        ctl_cal_fail    : in     vl_logic;
        ctl_cal_req     : out    vl_logic;
        ctl_init_req    : out    vl_logic;
        ctl_mem_clk_disable: out    vl_logic_vector;
        ctl_cal_byte_lane_sel_n: out    vl_logic_vector;
        cfg_type        : in     vl_logic_vector;
        cfg_interface_width: in     vl_logic_vector;
        cfg_burst_length: in     vl_logic_vector;
        cfg_device_width: in     vl_logic_vector;
        cfg_output_regd : in     vl_logic_vector;
        cfg_addr_order  : in     vl_logic_vector;
        cfg_col_addr_width: in     vl_logic_vector;
        cfg_row_addr_width: in     vl_logic_vector;
        cfg_bank_addr_width: in     vl_logic_vector;
        cfg_cs_addr_width: in     vl_logic_vector;
        cfg_cas_wr_lat  : in     vl_logic_vector;
        cfg_add_lat     : in     vl_logic_vector;
        cfg_tcl         : in     vl_logic_vector;
        cfg_trrd        : in     vl_logic_vector;
        cfg_tfaw        : in     vl_logic_vector;
        cfg_trfc        : in     vl_logic_vector;
        cfg_trefi       : in     vl_logic_vector;
        cfg_trcd        : in     vl_logic_vector;
        cfg_trp         : in     vl_logic_vector;
        cfg_twr         : in     vl_logic_vector;
        cfg_twtr        : in     vl_logic_vector;
        cfg_trtp        : in     vl_logic_vector;
        cfg_tras        : in     vl_logic_vector;
        cfg_trc         : in     vl_logic_vector;
        cfg_tccd        : in     vl_logic_vector;
        cfg_auto_pd_cycles: in     vl_logic_vector;
        cfg_self_rfsh_exit_cycles: in     vl_logic_vector;
        cfg_pdn_exit_cycles: in     vl_logic_vector;
        cfg_power_saving_exit_cycles: in     vl_logic_vector;
        cfg_mem_clk_entry_cycles: in     vl_logic_vector;
        cfg_tmrd        : in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_rdwr: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_pch: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_act: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_rd: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_rd_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_wr: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_wr_bc: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_wr_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_to_pch: in     vl_logic_vector;
        cfg_extra_ctl_clk_rd_ap_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_wr: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_wr_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_rd: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_rd_bc: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_rd_diff_chip: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_to_pch: in     vl_logic_vector;
        cfg_extra_ctl_clk_wr_ap_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_pch_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_pch_all_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_act_to_act_diff_bank: in     vl_logic_vector;
        cfg_extra_ctl_clk_four_act_to_act: in     vl_logic_vector;
        cfg_extra_ctl_clk_arf_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_pdn_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_srf_to_valid: in     vl_logic_vector;
        cfg_extra_ctl_clk_srf_to_zq_cal: in     vl_logic_vector;
        cfg_extra_ctl_clk_arf_period: in     vl_logic_vector;
        cfg_extra_ctl_clk_pdn_period: in     vl_logic_vector;
        cfg_reorder_data: in     vl_logic_vector;
        cfg_starve_limit: in     vl_logic_vector;
        cfg_user_rfsh   : in     vl_logic_vector;
        cfg_regdimm_enable: in     vl_logic_vector;
        cfg_enable_burst_interrupt: in     vl_logic_vector;
        cfg_enable_burst_terminate: in     vl_logic_vector;
        cfg_enable_ecc  : in     vl_logic_vector;
        cfg_enable_auto_corr: in     vl_logic_vector;
        cfg_enable_ecc_code_overwrites: in     vl_logic_vector;
        cfg_enable_no_dm: in     vl_logic_vector;
        cfg_gen_sbe     : in     vl_logic_vector;
        cfg_gen_dbe     : in     vl_logic_vector;
        cfg_enable_intr : in     vl_logic_vector;
        cfg_mask_sbe_intr: in     vl_logic_vector;
        cfg_mask_dbe_intr: in     vl_logic_vector;
        cfg_mask_corr_dropped_intr: in     vl_logic_vector;
        cfg_clr_intr    : in     vl_logic_vector;
        cfg_write_odt_chip: in     vl_logic_vector;
        cfg_read_odt_chip: in     vl_logic_vector;
        ecc_interrupt   : out    vl_logic;
        sts_sbe_error   : out    vl_logic_vector;
        sts_dbe_error   : out    vl_logic_vector;
        sts_corr_dropped: out    vl_logic_vector;
        sts_sbe_count   : out    vl_logic_vector;
        sts_dbe_count   : out    vl_logic_vector;
        sts_corr_dropped_count: out    vl_logic_vector;
        sts_err_addr    : out    vl_logic_vector;
        sts_corr_dropped_addr: out    vl_logic_vector;
        cfg_cal_req     : in     vl_logic;
        sts_cal_fail    : out    vl_logic;
        sts_cal_success : out    vl_logic;
        cfg_enable_dqs_tracking: in     vl_logic;
        afi_ctl_refresh_done: out    vl_logic_vector;
        afi_seq_busy    : in     vl_logic_vector;
        afi_ctl_long_idle: out    vl_logic_vector;
        tbp_empty       : out    vl_logic;
        cmd_gen_busy    : out    vl_logic;
        sideband_in_refresh: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_LOCAL_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_IF_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_BA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CKE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CLK_PAIR_COUNT : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_ODT_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of \CFG_OUTPUT_REGD\ : constant is 1;
    attribute mti_svvh_generic_type of CFG_CTL_TBP_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_LPDDR2_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_REORDERING_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_MULTIPLES_16_24_40_72 : constant is 1;
    attribute mti_svvh_generic_type of CFG_WRBUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_RDBUFFER_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MAX_PENDING_RD_CMD : constant is 1;
    attribute mti_svvh_generic_type of CFG_MAX_PENDING_WR_CMD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_INTERFACE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_BURST_LENGTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_DEVICE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_OUTPUT_REGD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ADDR_ORDER : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_COL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ROW_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_BANK_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_CS_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_CAS_WR_LAT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ADD_LAT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TCL : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRRD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TFAW : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRFC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TREFI : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRCD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TWR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TWTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRTP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRAS : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TRC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TCCD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TMRD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_SELF_RFSH_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_PDN_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_AUTO_PD_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_POWER_SAVING_EXIT_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MEM_CLK_ENTRY_CYCLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_RDWR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_PCH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_RD_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_BC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_WR_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_TO_PCH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_RD_AP_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_WR_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_BC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_RD_DIFF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_TO_PCH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_WR_AP_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PCH_ALL_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ACT_TO_ACT_DIFF_BANK : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_FOUR_ACT_TO_ACT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_VALID : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_SRF_TO_ZQ_CAL : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_ARF_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_EXTRA_CTL_CLK_PDN_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_REORDER_DATA : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_STARVE_LIMIT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_USER_RFSH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_SELF_RFSH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_REGDIMM_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_BURST_INTERRUPT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_BURST_TERMINATE : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_CMD_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_WDATA_PATH_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_ECC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_AUTO_CORR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_GEN_SBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_GEN_DBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MASK_SBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MASK_DBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MASK_CORR_DROPPED_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_CLR_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_ECC_CODE_OVERWRITES : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_NO_DM : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_DECODER_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_WRITE_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_READ_ODT_CHIP : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_SBE_ERROR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_DBE_ERROR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_CORR_DROP_ERROR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_SBE_COUNT : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_DBE_COUNT : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_CORR_DROP_COUNT : constant is 1;
    attribute mti_svvh_generic_type of CFG_WLAT_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_RRANK_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_WRANK_BUS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_USE_SHADOW_REGS : constant is 1;
    attribute mti_svvh_generic_type of CFG_RDATA_RETURN_MODE : constant is 1;
    attribute mti_svvh_generic_type of CFG_ERRCMD_FIFO_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_BURST_MERGE : constant is 1;
end alt_mem_ddrx_controller;
