library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_tbp is
    generic(
        CFG_CTL_TBP_NUM : integer := 4;
        CFG_CTL_SHADOW_TBP_NUM: integer := 4;
        CFG_ENABLE_SHADOW_TBP: integer := 0;
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_CTL_ARBITER_TYPE: string  := "ROWCOL";
        CFG_MEM_IF_CHIP : integer := 1;
        CFG_MEM_IF_CS_WIDTH: integer := 1;
        CFG_MEM_IF_BA_WIDTH: integer := 3;
        CFG_MEM_IF_ROW_WIDTH: integer := 13;
        CFG_MEM_IF_COL_WIDTH: integer := 10;
        CFG_LOCAL_ID_WIDTH: integer := 8;
        CFG_INT_SIZE_WIDTH: integer := 4;
        CFG_DATA_ID_WIDTH: integer := 10;
        CFG_REG_REQ     : integer := 0;
        CFG_REG_GRANT   : integer := 0;
        CFG_DATA_REORDERING_TYPE: string  := "INTER_BANK";
        CFG_DISABLE_READ_REODERING: integer := 0;
        CFG_DISABLE_PRIORITY: integer := 0;
        CFG_PORT_WIDTH_REORDER_DATA: integer := 1;
        CFG_PORT_WIDTH_STARVE_LIMIT: integer := 6;
        CFG_PORT_WIDTH_TYPE: integer := 3;
        T_PARAM_ACT_TO_RDWR_WIDTH: integer := 4;
        T_PARAM_ACT_TO_ACT_WIDTH: integer := 4;
        T_PARAM_ACT_TO_PCH_WIDTH: integer := 4;
        T_PARAM_RD_TO_PCH_WIDTH: integer := 4;
        T_PARAM_WR_TO_PCH_WIDTH: integer := 4;
        T_PARAM_PCH_TO_VALID_WIDTH: integer := 4;
        T_PARAM_RD_AP_TO_VALID_WIDTH: integer := 4;
        T_PARAM_WR_AP_TO_VALID_WIDTH: integer := 4
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        tbp_full        : out    vl_logic;
        tbp_empty       : out    vl_logic;
        cmd_gen_load    : in     vl_logic;
        cmd_gen_waiting_to_load: in     vl_logic;
        cmd_gen_chipsel : in     vl_logic_vector;
        cmd_gen_bank    : in     vl_logic_vector;
        cmd_gen_row     : in     vl_logic_vector;
        cmd_gen_col     : in     vl_logic_vector;
        cmd_gen_write   : in     vl_logic;
        cmd_gen_read    : in     vl_logic;
        cmd_gen_size    : in     vl_logic_vector;
        cmd_gen_localid : in     vl_logic_vector;
        cmd_gen_dataid  : in     vl_logic_vector;
        cmd_gen_priority: in     vl_logic;
        cmd_gen_rmw_correct: in     vl_logic;
        cmd_gen_rmw_partial: in     vl_logic;
        cmd_gen_autopch : in     vl_logic;
        cmd_gen_complete: in     vl_logic;
        cmd_gen_same_chipsel_addr: in     vl_logic_vector;
        cmd_gen_same_bank_addr: in     vl_logic_vector;
        cmd_gen_same_row_addr: in     vl_logic_vector;
        cmd_gen_same_col_addr: in     vl_logic_vector;
        cmd_gen_same_read_cmd: in     vl_logic_vector;
        cmd_gen_same_write_cmd: in     vl_logic_vector;
        cmd_gen_same_shadow_chipsel_addr: in     vl_logic_vector;
        cmd_gen_same_shadow_bank_addr: in     vl_logic_vector;
        cmd_gen_same_shadow_row_addr: in     vl_logic_vector;
        row_req         : out    vl_logic_vector;
        act_req         : out    vl_logic_vector;
        pch_req         : out    vl_logic_vector;
        row_grant       : in     vl_logic_vector;
        act_grant       : in     vl_logic_vector;
        pch_grant       : in     vl_logic_vector;
        col_req         : out    vl_logic_vector;
        rd_req          : out    vl_logic_vector;
        wr_req          : out    vl_logic_vector;
        col_grant       : in     vl_logic_vector;
        rd_grant        : in     vl_logic_vector;
        wr_grant        : in     vl_logic_vector;
        log2_row_grant  : in     vl_logic_vector;
        log2_col_grant  : in     vl_logic_vector;
        log2_act_grant  : in     vl_logic_vector;
        log2_pch_grant  : in     vl_logic_vector;
        log2_rd_grant   : in     vl_logic_vector;
        log2_wr_grant   : in     vl_logic_vector;
        or_row_grant    : in     vl_logic;
        or_col_grant    : in     vl_logic;
        tbp_read        : out    vl_logic_vector;
        tbp_write       : out    vl_logic_vector;
        tbp_precharge   : out    vl_logic_vector;
        tbp_activate    : out    vl_logic_vector;
        tbp_chipsel     : out    vl_logic_vector;
        tbp_bank        : out    vl_logic_vector;
        tbp_row         : out    vl_logic_vector;
        tbp_col         : out    vl_logic_vector;
        tbp_shadow_chipsel: out    vl_logic_vector;
        tbp_shadow_bank : out    vl_logic_vector;
        tbp_shadow_row  : out    vl_logic_vector;
        tbp_size        : out    vl_logic_vector;
        tbp_localid     : out    vl_logic_vector;
        tbp_dataid      : out    vl_logic_vector;
        tbp_ap          : out    vl_logic_vector;
        tbp_burst_chop  : out    vl_logic_vector;
        tbp_age         : out    vl_logic_vector;
        tbp_priority    : out    vl_logic_vector;
        tbp_rmw_correct : out    vl_logic_vector;
        tbp_rmw_partial : out    vl_logic_vector;
        sb_tbp_precharge_all: in     vl_logic_vector;
        sb_do_precharge_all: in     vl_logic_vector;
        t_param_act_to_rdwr: in     vl_logic_vector;
        t_param_act_to_act: in     vl_logic_vector;
        t_param_act_to_pch: in     vl_logic_vector;
        t_param_rd_to_pch: in     vl_logic_vector;
        t_param_wr_to_pch: in     vl_logic_vector;
        t_param_pch_to_valid: in     vl_logic_vector;
        t_param_rd_ap_to_valid: in     vl_logic_vector;
        t_param_wr_ap_to_valid: in     vl_logic_vector;
        tbp_bank_closed : out    vl_logic_vector;
        tbp_timer_ready : out    vl_logic_vector;
        tbp_load        : out    vl_logic_vector;
        data_complete   : in     vl_logic_vector;
        data_rmw_complete: in     vl_logic;
        data_rmw_fetch  : out    vl_logic;
        cfg_reorder_data: in     vl_logic_vector;
        cfg_starve_limit: in     vl_logic_vector;
        cfg_type        : in     vl_logic_vector;
        cfg_enable_ecc  : in     vl_logic;
        cfg_enable_no_dm: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_CTL_TBP_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_CTL_SHADOW_TBP_NUM : constant is 1;
    attribute mti_svvh_generic_type of CFG_ENABLE_SHADOW_TBP : constant is 1;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_CTL_ARBITER_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CHIP : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_BA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_ROW_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_COL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_INT_SIZE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_ID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_REG_REQ : constant is 1;
    attribute mti_svvh_generic_type of CFG_REG_GRANT : constant is 1;
    attribute mti_svvh_generic_type of CFG_DATA_REORDERING_TYPE : constant is 1;
    attribute mti_svvh_generic_type of CFG_DISABLE_READ_REODERING : constant is 1;
    attribute mti_svvh_generic_type of CFG_DISABLE_PRIORITY : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_REORDER_DATA : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_STARVE_LIMIT : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_TYPE : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_RDWR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_ACT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_ACT_TO_PCH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_TO_PCH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_TO_PCH_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_PCH_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_RD_AP_TO_VALID_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of T_PARAM_WR_AP_TO_VALID_WIDTH : constant is 1;
end alt_mem_ddrx_tbp;
