library verilog;
use verilog.vl_types.all;
entity altera_conduit_bfm_0004 is
    port(
        sig_export      : out    vl_logic_vector(3 downto 0)
    );
end altera_conduit_bfm_0004;
