library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_tb is
end DE4_QSYS_tb;
