// DE4_QSYS.v

// Generated using ACDS version 13.0sp1 232 at 2015.07.12.17:21:47

`timescale 1 ps / 1 ps
module DE4_QSYS (
		input  wire        clk_clk,                                   //                     clk.clk
		input  wire        reset_reset_n,                             //                   reset.reset_n
		output wire [13:0] memory_mem_a,                              //                  memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                        .mem_ba
		output wire [1:0]  memory_mem_ck,                             //                        .mem_ck
		output wire [1:0]  memory_mem_ck_n,                           //                        .mem_ck_n
		output wire [0:0]  memory_mem_cke,                            //                        .mem_cke
		output wire [0:0]  memory_mem_cs_n,                           //                        .mem_cs_n
		output wire [7:0]  memory_mem_dm,                             //                        .mem_dm
		output wire [0:0]  memory_mem_ras_n,                          //                        .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                          //                        .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                           //                        .mem_we_n
		inout  wire [63:0] memory_mem_dq,                             //                        .mem_dq
		inout  wire [7:0]  memory_mem_dqs,                            //                        .mem_dqs
		inout  wire [7:0]  memory_mem_dqs_n,                          //                        .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                            //                        .mem_odt
		input  wire        oct_rdn,                                   //                     oct.rdn
		input  wire        oct_rup,                                   //                        .rup
		output wire        mem_if_ddr2_emif_status_local_init_done,   // mem_if_ddr2_emif_status.local_init_done
		output wire        mem_if_ddr2_emif_status_local_cal_success, //                        .local_cal_success
		output wire        mem_if_ddr2_emif_status_local_cal_fail,    //                        .local_cal_fail
		output wire [7:0]  led_export,                                //                     led.export
		input  wire [3:0]  button_export,                             //                  button.export
		output wire        ddr2_i2c_scl_export,                       //            ddr2_i2c_scl.export
		inout  wire        ddr2_i2c_sda_export                        //            ddr2_i2c_sda.export
	);

	wire          mem_if_ddr2_emif_afi_clk_clk;                                                                        // mem_if_ddr2_emif:afi_clk -> [addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, addr_router_005:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_demux_005:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_004:clk, crosser:in_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:in_clk, crosser_005:in_clk, crosser_006:in_clk, crosser_007:in_clk, crosser_008:out_clk, crosser_009:out_clk, crosser_010:out_clk, crosser_011:out_clk, crosser_012:out_clk, crosser_013:out_clk, dma:clk, dma_control_port_slave_translator:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dma_read_master_translator:clk, dma_read_master_translator_avalon_universal_master_0_agent:clk, dma_write_master_translator:clk, dma_write_master_translator_avalon_universal_master_0_agent:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, limiter_002:clk, mem_if_ddr2_emif_avl_translator:clk, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:clk, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, mm_clock_crossing_bridge_io:m0_clk, mm_clock_crossing_bridge_io_m0_translator:clk, mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:clk, nios2_qsys:clk, nios2_qsys_data_master_translator:clk, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_instruction_master_translator:clk, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_jtag_debug_module_translator:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory:clk, onchip_memory_s1_translator:clk, onchip_memory_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ppl_mem_reader:clk, ppl_mem_reader_avalon_master_translator:clk, ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_005:clk, rst_controller:clk, rst_controller_002:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, wrapper_0:clk, wrapper_0_s0_translator:clk, wrapper_0_s0_translator_avalon_universal_slave_0_agent:clk, wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire          wrapper_0_control_fixed_location;                                                                    // wrapper_0:coe_control_fixed_location -> ppl_mem_reader:coe_control_fixed_location
	wire   [31:0] wrapper_0_control_read_base;                                                                         // wrapper_0:coe_control_read_base -> ppl_mem_reader:coe_control_read_base
	wire          ppl_mem_reader_control_early_done;                                                                   // ppl_mem_reader:coe_control_early_done -> wrapper_0:coe_control_early_done
	wire          ppl_mem_reader_control_done;                                                                         // ppl_mem_reader:coe_control_done -> wrapper_0:coe_control_done
	wire   [31:0] wrapper_0_control_read_length;                                                                       // wrapper_0:coe_control_read_length -> ppl_mem_reader:coe_control_read_length
	wire          wrapper_0_control_go;                                                                                // wrapper_0:coe_control_go -> ppl_mem_reader:coe_control_go
	wire          wrapper_0_user_read_buffer;                                                                          // wrapper_0:coe_user_read_buffer -> ppl_mem_reader:coe_user_read_buffer
	wire   [31:0] ppl_mem_reader_user_buffer_data;                                                                     // ppl_mem_reader:coe_user_buffer_data -> wrapper_0:coe_user_buffer_data
	wire          ppl_mem_reader_user_data_available;                                                                  // ppl_mem_reader:coe_user_data_available -> wrapper_0:coe_user_data_available
	wire          nios2_qsys_instruction_master_waitrequest;                                                           // nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	wire   [30:0] nios2_qsys_instruction_master_address;                                                               // nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	wire          nios2_qsys_instruction_master_read;                                                                  // nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	wire   [31:0] nios2_qsys_instruction_master_readdata;                                                              // nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	wire          nios2_qsys_instruction_master_readdatavalid;                                                         // nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	wire    [3:0] nios2_qsys_data_master_burstcount;                                                                   // nios2_qsys:d_burstcount -> nios2_qsys_data_master_translator:av_burstcount
	wire          nios2_qsys_data_master_waitrequest;                                                                  // nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	wire   [31:0] nios2_qsys_data_master_writedata;                                                                    // nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	wire   [30:0] nios2_qsys_data_master_address;                                                                      // nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	wire          nios2_qsys_data_master_write;                                                                        // nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	wire          nios2_qsys_data_master_read;                                                                         // nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	wire   [31:0] nios2_qsys_data_master_readdata;                                                                     // nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	wire          nios2_qsys_data_master_debugaccess;                                                                  // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	wire          nios2_qsys_data_master_readdatavalid;                                                                // nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	wire    [3:0] nios2_qsys_data_master_byteenable;                                                                   // nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	wire          dma_read_master_burstcount;                                                                          // dma:read_burstcount -> dma_read_master_translator:av_burstcount
	wire          dma_read_master_waitrequest;                                                                         // dma_read_master_translator:av_waitrequest -> dma:read_waitrequest
	wire   [29:0] dma_read_master_address;                                                                             // dma:read_address -> dma_read_master_translator:av_address
	wire          dma_read_master_chipselect;                                                                          // dma:read_chipselect -> dma_read_master_translator:av_chipselect
	wire          dma_read_master_read;                                                                                // dma:read_read_n -> dma_read_master_translator:av_read
	wire   [15:0] dma_read_master_readdata;                                                                            // dma_read_master_translator:av_readdata -> dma:read_readdata
	wire          dma_read_master_readdatavalid;                                                                       // dma_read_master_translator:av_readdatavalid -> dma:read_readdatavalid
	wire          dma_write_master_burstcount;                                                                         // dma:write_burstcount -> dma_write_master_translator:av_burstcount
	wire          dma_write_master_waitrequest;                                                                        // dma_write_master_translator:av_waitrequest -> dma:write_waitrequest
	wire   [15:0] dma_write_master_writedata;                                                                          // dma:write_writedata -> dma_write_master_translator:av_writedata
	wire   [29:0] dma_write_master_address;                                                                            // dma:write_address -> dma_write_master_translator:av_address
	wire          dma_write_master_chipselect;                                                                         // dma:write_chipselect -> dma_write_master_translator:av_chipselect
	wire          dma_write_master_write;                                                                              // dma:write_write_n -> dma_write_master_translator:av_write
	wire    [1:0] dma_write_master_byteenable;                                                                         // dma:write_byteenable -> dma_write_master_translator:av_byteenable
	wire          ppl_mem_reader_avalon_master_waitrequest;                                                            // ppl_mem_reader_avalon_master_translator:av_waitrequest -> ppl_mem_reader:master_waitrequest
	wire   [31:0] ppl_mem_reader_avalon_master_address;                                                                // ppl_mem_reader:master_address -> ppl_mem_reader_avalon_master_translator:av_address
	wire          ppl_mem_reader_avalon_master_read;                                                                   // ppl_mem_reader:master_read -> ppl_mem_reader_avalon_master_translator:av_read
	wire   [31:0] ppl_mem_reader_avalon_master_readdata;                                                               // ppl_mem_reader_avalon_master_translator:av_readdata -> ppl_mem_reader:master_readdata
	wire          ppl_mem_reader_avalon_master_readdatavalid;                                                          // ppl_mem_reader_avalon_master_translator:av_readdatavalid -> ppl_mem_reader:master_readdatavalid
	wire    [3:0] ppl_mem_reader_avalon_master_byteenable;                                                             // ppl_mem_reader:master_byteenable -> ppl_mem_reader_avalon_master_translator:av_byteenable
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                             // nios2_qsys:jtag_debug_module_waitrequest -> nios2_qsys_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                               // nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire    [8:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address;                                 // nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write;                                   // nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read;                                    // nios2_qsys_jtag_debug_module_translator:av_read -> nios2_qsys:jtag_debug_module_read
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                // nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	wire          nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                             // nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire    [3:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                              // nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_writedata;                                           // onchip_memory_s1_translator:av_writedata -> onchip_memory:writedata
	wire   [14:0] onchip_memory_s1_translator_avalon_anti_slave_0_address;                                             // onchip_memory_s1_translator:av_address -> onchip_memory:address
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_chipselect;                                          // onchip_memory_s1_translator:av_chipselect -> onchip_memory:chipselect
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_clken;                                               // onchip_memory_s1_translator:av_clken -> onchip_memory:clken
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_write;                                               // onchip_memory_s1_translator:av_write -> onchip_memory:write
	wire   [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_readdata;                                            // onchip_memory:readdata -> onchip_memory_s1_translator:av_readdata
	wire    [3:0] onchip_memory_s1_translator_avalon_anti_slave_0_byteenable;                                          // onchip_memory_s1_translator:av_byteenable -> onchip_memory:byteenable
	wire   [30:0] dma_control_port_slave_translator_avalon_anti_slave_0_writedata;                                     // dma_control_port_slave_translator:av_writedata -> dma:dma_ctl_writedata
	wire    [2:0] dma_control_port_slave_translator_avalon_anti_slave_0_address;                                       // dma_control_port_slave_translator:av_address -> dma:dma_ctl_address
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                    // dma_control_port_slave_translator:av_chipselect -> dma:dma_ctl_chipselect
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_write;                                         // dma_control_port_slave_translator:av_write -> dma:dma_ctl_write_n
	wire   [30:0] dma_control_port_slave_translator_avalon_anti_slave_0_readdata;                                      // dma:dma_ctl_readdata -> dma_control_port_slave_translator:av_readdata
	wire   [31:0] wrapper_0_s0_translator_avalon_anti_slave_0_writedata;                                               // wrapper_0_s0_translator:av_writedata -> wrapper_0:avs_s0_writedata
	wire    [1:0] wrapper_0_s0_translator_avalon_anti_slave_0_address;                                                 // wrapper_0_s0_translator:av_address -> wrapper_0:avs_s0_address
	wire          wrapper_0_s0_translator_avalon_anti_slave_0_write;                                                   // wrapper_0_s0_translator:av_write -> wrapper_0:avs_s0_write
	wire          wrapper_0_s0_translator_avalon_anti_slave_0_read;                                                    // wrapper_0_s0_translator:av_read -> wrapper_0:avs_s0_read
	wire   [31:0] wrapper_0_s0_translator_avalon_anti_slave_0_readdata;                                                // wrapper_0:avs_s0_readdata -> wrapper_0_s0_translator:av_readdata
	wire          wrapper_0_s0_translator_avalon_anti_slave_0_readdatavalid;                                           // wrapper_0:avs_s0_readdatavalid -> wrapper_0_s0_translator:av_readdatavalid
	wire          mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_waitrequest;                                     // mem_if_ddr2_emif:avl_ready -> mem_if_ddr2_emif_avl_translator:av_waitrequest
	wire    [2:0] mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_burstcount;                                      // mem_if_ddr2_emif_avl_translator:av_burstcount -> mem_if_ddr2_emif:avl_size
	wire  [255:0] mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_writedata;                                       // mem_if_ddr2_emif_avl_translator:av_writedata -> mem_if_ddr2_emif:avl_wdata
	wire   [24:0] mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_address;                                         // mem_if_ddr2_emif_avl_translator:av_address -> mem_if_ddr2_emif:avl_addr
	wire          mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_write;                                           // mem_if_ddr2_emif_avl_translator:av_write -> mem_if_ddr2_emif:avl_write_req
	wire          mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_beginbursttransfer;                              // mem_if_ddr2_emif_avl_translator:av_beginbursttransfer -> mem_if_ddr2_emif:avl_burstbegin
	wire          mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_read;                                            // mem_if_ddr2_emif_avl_translator:av_read -> mem_if_ddr2_emif:avl_read_req
	wire  [255:0] mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdata;                                        // mem_if_ddr2_emif:avl_rdata -> mem_if_ddr2_emif_avl_translator:av_readdata
	wire          mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdatavalid;                                   // mem_if_ddr2_emif:avl_rdata_valid -> mem_if_ddr2_emif_avl_translator:av_readdatavalid
	wire   [31:0] mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_byteenable;                                      // mem_if_ddr2_emif_avl_translator:av_byteenable -> mem_if_ddr2_emif:avl_be
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                              // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                  // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                               // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                    // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                     // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                 // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_waitrequest;                           // mm_clock_crossing_bridge_io:s0_waitrequest -> mm_clock_crossing_bridge_io_s0_translator:av_waitrequest
	wire    [0:0] mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_burstcount;                            // mm_clock_crossing_bridge_io_s0_translator:av_burstcount -> mm_clock_crossing_bridge_io:s0_burstcount
	wire   [31:0] mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_writedata;                             // mm_clock_crossing_bridge_io_s0_translator:av_writedata -> mm_clock_crossing_bridge_io:s0_writedata
	wire    [9:0] mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_address;                               // mm_clock_crossing_bridge_io_s0_translator:av_address -> mm_clock_crossing_bridge_io:s0_address
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_write;                                 // mm_clock_crossing_bridge_io_s0_translator:av_write -> mm_clock_crossing_bridge_io:s0_write
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_read;                                  // mm_clock_crossing_bridge_io_s0_translator:av_read -> mm_clock_crossing_bridge_io:s0_read
	wire   [31:0] mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdata;                              // mm_clock_crossing_bridge_io:s0_readdata -> mm_clock_crossing_bridge_io_s0_translator:av_readdata
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_debugaccess;                           // mm_clock_crossing_bridge_io_s0_translator:av_debugaccess -> mm_clock_crossing_bridge_io:s0_debugaccess
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdatavalid;                         // mm_clock_crossing_bridge_io:s0_readdatavalid -> mm_clock_crossing_bridge_io_s0_translator:av_readdatavalid
	wire    [3:0] mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_byteenable;                            // mm_clock_crossing_bridge_io_s0_translator:av_byteenable -> mm_clock_crossing_bridge_io:s0_byteenable
	wire    [0:0] mm_clock_crossing_bridge_io_m0_burstcount;                                                           // mm_clock_crossing_bridge_io:m0_burstcount -> mm_clock_crossing_bridge_io_m0_translator:av_burstcount
	wire          mm_clock_crossing_bridge_io_m0_waitrequest;                                                          // mm_clock_crossing_bridge_io_m0_translator:av_waitrequest -> mm_clock_crossing_bridge_io:m0_waitrequest
	wire    [9:0] mm_clock_crossing_bridge_io_m0_address;                                                              // mm_clock_crossing_bridge_io:m0_address -> mm_clock_crossing_bridge_io_m0_translator:av_address
	wire   [31:0] mm_clock_crossing_bridge_io_m0_writedata;                                                            // mm_clock_crossing_bridge_io:m0_writedata -> mm_clock_crossing_bridge_io_m0_translator:av_writedata
	wire          mm_clock_crossing_bridge_io_m0_write;                                                                // mm_clock_crossing_bridge_io:m0_write -> mm_clock_crossing_bridge_io_m0_translator:av_write
	wire          mm_clock_crossing_bridge_io_m0_read;                                                                 // mm_clock_crossing_bridge_io:m0_read -> mm_clock_crossing_bridge_io_m0_translator:av_read
	wire   [31:0] mm_clock_crossing_bridge_io_m0_readdata;                                                             // mm_clock_crossing_bridge_io_m0_translator:av_readdata -> mm_clock_crossing_bridge_io:m0_readdata
	wire          mm_clock_crossing_bridge_io_m0_debugaccess;                                                          // mm_clock_crossing_bridge_io:m0_debugaccess -> mm_clock_crossing_bridge_io_m0_translator:av_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_io_m0_byteenable;                                                           // mm_clock_crossing_bridge_io:m0_byteenable -> mm_clock_crossing_bridge_io_m0_translator:av_byteenable
	wire          mm_clock_crossing_bridge_io_m0_readdatavalid;                                                        // mm_clock_crossing_bridge_io_m0_translator:av_readdatavalid -> mm_clock_crossing_bridge_io:m0_readdatavalid
	wire    [1:0] button_s1_translator_avalon_anti_slave_0_address;                                                    // button_s1_translator:av_address -> button:address
	wire   [31:0] button_s1_translator_avalon_anti_slave_0_readdata;                                                   // button:readdata -> button_s1_translator:av_readdata
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                                                     // led_s1_translator:av_writedata -> led:writedata
	wire    [1:0] led_s1_translator_avalon_anti_slave_0_address;                                                       // led_s1_translator:av_address -> led:address
	wire          led_s1_translator_avalon_anti_slave_0_chipselect;                                                    // led_s1_translator:av_chipselect -> led:chipselect
	wire          led_s1_translator_avalon_anti_slave_0_write;                                                         // led_s1_translator:av_write -> led:write_n
	wire   [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                                                      // led:readdata -> led_s1_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                   // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                     // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                                  // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                       // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                    // timer:readdata -> timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                          // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                         // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                            // ddr2_i2c_scl_s1_translator:av_writedata -> ddr2_i2c_scl:writedata
	wire    [1:0] ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_address;                                              // ddr2_i2c_scl_s1_translator:av_address -> ddr2_i2c_scl:address
	wire          ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                           // ddr2_i2c_scl_s1_translator:av_chipselect -> ddr2_i2c_scl:chipselect
	wire          ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                // ddr2_i2c_scl_s1_translator:av_write -> ddr2_i2c_scl:write_n
	wire   [31:0] ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                             // ddr2_i2c_scl:readdata -> ddr2_i2c_scl_s1_translator:av_readdata
	wire   [31:0] ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                            // ddr2_i2c_sda_s1_translator:av_writedata -> ddr2_i2c_sda:writedata
	wire    [1:0] ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_address;                                              // ddr2_i2c_sda_s1_translator:av_address -> ddr2_i2c_sda:address
	wire          ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                           // ddr2_i2c_sda_s1_translator:av_chipselect -> ddr2_i2c_sda:chipselect
	wire          ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_write;                                                // ddr2_i2c_sda_s1_translator:av_write -> ddr2_i2c_sda:write_n
	wire   [31:0] ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                             // ddr2_i2c_sda:readdata -> ddr2_i2c_sda_s1_translator:av_readdata
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest;                      // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount;                       // nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata;                        // nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_address;                          // nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock;                             // nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_write;                            // nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_read;                             // nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata;                         // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess;                      // nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable;                       // nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid;                    // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest;                             // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	wire    [5:0] nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount;                              // nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_writedata;                               // nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_address;                                 // nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_lock;                                    // nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_write;                                   // nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_read;                                    // nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_readdata;                                // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess;                             // nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable;                              // nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid;                           // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	wire          dma_read_master_translator_avalon_universal_master_0_waitrequest;                                    // dma_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_read_master_translator:uav_waitrequest
	wire    [1:0] dma_read_master_translator_avalon_universal_master_0_burstcount;                                     // dma_read_master_translator:uav_burstcount -> dma_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] dma_read_master_translator_avalon_universal_master_0_writedata;                                      // dma_read_master_translator:uav_writedata -> dma_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_address;                                        // dma_read_master_translator:uav_address -> dma_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_read_master_translator_avalon_universal_master_0_lock;                                           // dma_read_master_translator:uav_lock -> dma_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_read_master_translator_avalon_universal_master_0_write;                                          // dma_read_master_translator:uav_write -> dma_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_read_master_translator_avalon_universal_master_0_read;                                           // dma_read_master_translator:uav_read -> dma_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] dma_read_master_translator_avalon_universal_master_0_readdata;                                       // dma_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_read_master_translator:uav_readdata
	wire          dma_read_master_translator_avalon_universal_master_0_debugaccess;                                    // dma_read_master_translator:uav_debugaccess -> dma_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] dma_read_master_translator_avalon_universal_master_0_byteenable;                                     // dma_read_master_translator:uav_byteenable -> dma_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_read_master_translator_avalon_universal_master_0_readdatavalid;                                  // dma_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_read_master_translator:uav_readdatavalid
	wire          dma_write_master_translator_avalon_universal_master_0_waitrequest;                                   // dma_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_write_master_translator:uav_waitrequest
	wire    [1:0] dma_write_master_translator_avalon_universal_master_0_burstcount;                                    // dma_write_master_translator:uav_burstcount -> dma_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] dma_write_master_translator_avalon_universal_master_0_writedata;                                     // dma_write_master_translator:uav_writedata -> dma_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_address;                                       // dma_write_master_translator:uav_address -> dma_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_write_master_translator_avalon_universal_master_0_lock;                                          // dma_write_master_translator:uav_lock -> dma_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_write_master_translator_avalon_universal_master_0_write;                                         // dma_write_master_translator:uav_write -> dma_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_write_master_translator_avalon_universal_master_0_read;                                          // dma_write_master_translator:uav_read -> dma_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] dma_write_master_translator_avalon_universal_master_0_readdata;                                      // dma_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_write_master_translator:uav_readdata
	wire          dma_write_master_translator_avalon_universal_master_0_debugaccess;                                   // dma_write_master_translator:uav_debugaccess -> dma_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] dma_write_master_translator_avalon_universal_master_0_byteenable;                                    // dma_write_master_translator:uav_byteenable -> dma_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_write_master_translator_avalon_universal_master_0_readdatavalid;                                 // dma_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_write_master_translator:uav_readdatavalid
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_waitrequest;                       // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> ppl_mem_reader_avalon_master_translator:uav_waitrequest
	wire    [2:0] ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_burstcount;                        // ppl_mem_reader_avalon_master_translator:uav_burstcount -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_writedata;                         // ppl_mem_reader_avalon_master_translator:uav_writedata -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_address;                           // ppl_mem_reader_avalon_master_translator:uav_address -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_lock;                              // ppl_mem_reader_avalon_master_translator:uav_lock -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_write;                             // ppl_mem_reader_avalon_master_translator:uav_write -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_read;                              // ppl_mem_reader_avalon_master_translator:uav_read -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_readdata;                          // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> ppl_mem_reader_avalon_master_translator:uav_readdata
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_debugaccess;                       // ppl_mem_reader_avalon_master_translator:uav_debugaccess -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_byteenable;                        // ppl_mem_reader_avalon_master_translator:uav_byteenable -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_readdatavalid;                     // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> ppl_mem_reader_avalon_master_translator:uav_readdatavalid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                 // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                     // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                  // nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [110:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [110:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // onchip_memory_s1_translator:uav_waitrequest -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_s1_translator:uav_writedata
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_s1_translator:uav_address
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_s1_translator:uav_write
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_s1_translator:uav_lock
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_s1_translator:uav_read
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // onchip_memory_s1_translator:uav_readdata -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // onchip_memory_s1_translator:uav_readdatavalid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_s1_translator:uav_byteenable
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [110:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [110:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // dma_control_port_slave_translator:uav_waitrequest -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_control_port_slave_translator:uav_writedata
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_control_port_slave_translator:uav_address
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_control_port_slave_translator:uav_write
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_control_port_slave_translator:uav_lock
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_control_port_slave_translator:uav_read
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // dma_control_port_slave_translator:uav_readdata -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // dma_control_port_slave_translator:uav_readdatavalid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_control_port_slave_translator:uav_byteenable
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [110:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [110:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // wrapper_0_s0_translator:uav_waitrequest -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> wrapper_0_s0_translator:uav_burstcount
	wire   [31:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> wrapper_0_s0_translator:uav_writedata
	wire   [31:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                                   // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> wrapper_0_s0_translator:uav_address
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                                     // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> wrapper_0_s0_translator:uav_write
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                      // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> wrapper_0_s0_translator:uav_lock
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                                      // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> wrapper_0_s0_translator:uav_read
	wire   [31:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // wrapper_0_s0_translator:uav_readdata -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // wrapper_0_s0_translator:uav_readdatavalid -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> wrapper_0_s0_translator:uav_debugaccess
	wire    [3:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // wrapper_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> wrapper_0_s0_translator:uav_byteenable
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [110:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                               // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [110:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // mem_if_ddr2_emif_avl_translator:uav_waitrequest -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [7:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> mem_if_ddr2_emif_avl_translator:uav_burstcount
	wire  [255:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_writedata;                         // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> mem_if_ddr2_emif_avl_translator:uav_writedata
	wire   [31:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_address;                           // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_address -> mem_if_ddr2_emif_avl_translator:uav_address
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_write;                             // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_write -> mem_if_ddr2_emif_avl_translator:uav_write
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_lock;                              // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_lock -> mem_if_ddr2_emif_avl_translator:uav_lock
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_read;                              // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_read -> mem_if_ddr2_emif_avl_translator:uav_read
	wire  [255:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                          // mem_if_ddr2_emif_avl_translator:uav_readdata -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // mem_if_ddr2_emif_avl_translator:uav_readdatavalid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mem_if_ddr2_emif_avl_translator:uav_debugaccess
	wire   [31:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> mem_if_ddr2_emif_avl_translator:uav_byteenable
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [362:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_data;                       // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [362:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [257:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [257:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [110:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [110:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // mm_clock_crossing_bridge_io_s0_translator:uav_waitrequest -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> mm_clock_crossing_bridge_io_s0_translator:uav_burstcount
	wire   [31:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata;               // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> mm_clock_crossing_bridge_io_s0_translator:uav_writedata
	wire   [31:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_address;                 // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_address -> mm_clock_crossing_bridge_io_s0_translator:uav_address
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_write;                   // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_write -> mm_clock_crossing_bridge_io_s0_translator:uav_write
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_lock;                    // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_lock -> mm_clock_crossing_bridge_io_s0_translator:uav_lock
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_read;                    // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_read -> mm_clock_crossing_bridge_io_s0_translator:uav_read
	wire   [31:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                // mm_clock_crossing_bridge_io_s0_translator:uav_readdata -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // mm_clock_crossing_bridge_io_s0_translator:uav_readdatavalid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mm_clock_crossing_bridge_io_s0_translator:uav_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> mm_clock_crossing_bridge_io_s0_translator:uav_byteenable
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [110:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data;             // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [110:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_waitrequest;                     // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> mm_clock_crossing_bridge_io_m0_translator:uav_waitrequest
	wire    [2:0] mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_burstcount;                      // mm_clock_crossing_bridge_io_m0_translator:uav_burstcount -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_writedata;                       // mm_clock_crossing_bridge_io_m0_translator:uav_writedata -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_address;                         // mm_clock_crossing_bridge_io_m0_translator:uav_address -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_address
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_lock;                            // mm_clock_crossing_bridge_io_m0_translator:uav_lock -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_write;                           // mm_clock_crossing_bridge_io_m0_translator:uav_write -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_write
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_read;                            // mm_clock_crossing_bridge_io_m0_translator:uav_read -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdata;                        // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_readdata -> mm_clock_crossing_bridge_io_m0_translator:uav_readdata
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_debugaccess;                     // mm_clock_crossing_bridge_io_m0_translator:uav_debugaccess -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_byteenable;                      // mm_clock_crossing_bridge_io_m0_translator:uav_byteenable -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdatavalid;                   // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> mm_clock_crossing_bridge_io_m0_translator:uav_readdatavalid
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // button_s1_translator:uav_waitrequest -> button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_s1_translator:uav_burstcount
	wire   [31:0] button_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_s1_translator:uav_writedata
	wire    [9:0] button_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // button_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_s1_translator:uav_address
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // button_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_s1_translator:uav_write
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_s1_translator:uav_lock
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // button_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_s1_translator:uav_read
	wire   [31:0] button_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // button_s1_translator:uav_readdata -> button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // button_s1_translator:uav_readdatavalid -> button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_s1_translator:uav_debugaccess
	wire    [3:0] button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_s1_translator:uav_byteenable
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] button_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                            // button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                             // button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                            // button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	wire    [9:0] led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	wire   [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	wire    [3:0] led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                               // led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                // led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                               // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire    [9:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                             // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                              // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                             // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [9:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // ddr2_i2c_scl_s1_translator:uav_waitrequest -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_i2c_scl_s1_translator:uav_burstcount
	wire   [31:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_i2c_scl_s1_translator:uav_writedata
	wire    [9:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_i2c_scl_s1_translator:uav_address
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_i2c_scl_s1_translator:uav_write
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_i2c_scl_s1_translator:uav_lock
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_i2c_scl_s1_translator:uav_read
	wire   [31:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // ddr2_i2c_scl_s1_translator:uav_readdata -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // ddr2_i2c_scl_s1_translator:uav_readdatavalid -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_i2c_scl_s1_translator:uav_debugaccess
	wire    [3:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_i2c_scl_s1_translator:uav_byteenable
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                      // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                       // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                      // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // ddr2_i2c_sda_s1_translator:uav_waitrequest -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_i2c_sda_s1_translator:uav_burstcount
	wire   [31:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_i2c_sda_s1_translator:uav_writedata
	wire    [9:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_i2c_sda_s1_translator:uav_address
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_i2c_sda_s1_translator:uav_write
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_i2c_sda_s1_translator:uav_lock
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_i2c_sda_s1_translator:uav_read
	wire   [31:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // ddr2_i2c_sda_s1_translator:uav_readdata -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // ddr2_i2c_sda_s1_translator:uav_readdatavalid -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_i2c_sda_s1_translator:uav_debugaccess
	wire    [3:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_i2c_sda_s1_translator:uav_byteenable
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [81:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [81:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                      // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                       // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                      // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;             // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                   // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;           // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [109:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                    // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                   // addr_router:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                    // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid;                          // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                  // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [109:0] nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data;                           // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready;                          // addr_router_001:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                           // dma_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_valid;                                 // dma_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                         // dma_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [91:0] dma_read_master_translator_avalon_universal_master_0_agent_cp_data;                                  // dma_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_ready;                                 // addr_router_002:sink_ready -> dma_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                          // dma_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_valid;                                // dma_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                        // dma_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [91:0] dma_write_master_translator_avalon_universal_master_0_agent_cp_data;                                 // dma_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_ready;                                // addr_router_003:sink_ready -> dma_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;              // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                    // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;            // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [109:0] ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                     // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router_004:sink_ready -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                     // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [109:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [109:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_001:sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [109:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_002:sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                     // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [109:0] wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                                      // wrapper_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_003:sink_ready -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_valid;                             // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [361:0] mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_data;                              // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_004:sink_ready -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [109:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_005:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_valid;                   // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [109:0] mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_data;                    // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;            // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_valid;                  // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;          // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire   [80:0] mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_data;                   // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router_005:sink_ready -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [80:0] button_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          button_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_007:sink_ready -> button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [80:0] led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_008:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [80:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_009:sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [80:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_010:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [80:0] ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_011:sink_ready -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [80:0] ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_012:sink_ready -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                               // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [109:0] addr_router_src_data;                                                                                // addr_router:src_data -> limiter:cmd_sink_data
	wire    [6:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                               // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                         // limiter:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                               // limiter:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                       // limiter:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [109:0] limiter_rsp_src_data;                                                                                // limiter:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [6:0] limiter_rsp_src_channel;                                                                             // limiter:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                               // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [109:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire    [6:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                           // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                     // limiter_001:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                           // limiter_001:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                   // limiter_001:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [109:0] limiter_001_rsp_src_data;                                                                            // limiter_001:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [6:0] limiter_001_rsp_src_channel;                                                                         // limiter_001:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                           // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_005_src_endofpacket;                                                                     // addr_router_005:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_005_src_valid;                                                                           // addr_router_005:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_005_src_startofpacket;                                                                   // addr_router_005:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [80:0] addr_router_005_src_data;                                                                            // addr_router_005:src_data -> limiter_002:cmd_sink_data
	wire    [5:0] addr_router_005_src_channel;                                                                         // addr_router_005:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_005_src_ready;                                                                           // limiter_002:cmd_sink_ready -> addr_router_005:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                     // limiter_002:rsp_src_endofpacket -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                           // limiter_002:rsp_src_valid -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                   // limiter_002:rsp_src_startofpacket -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [80:0] limiter_002_rsp_src_data;                                                                            // limiter_002:rsp_src_data -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_002_rsp_src_channel;                                                                         // limiter_002:rsp_src_channel -> mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                           // mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                   // burst_adapter:source0_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                         // burst_adapter:source0_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                 // burst_adapter:source0_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [109:0] burst_adapter_source0_data;                                                                          // burst_adapter:source0_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [6:0] burst_adapter_source0_channel;                                                                       // burst_adapter:source0_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                               // burst_adapter_001:source0_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                     // burst_adapter_001:source0_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                             // burst_adapter_001:source0_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [109:0] burst_adapter_001_source0_data;                                                                      // burst_adapter_001:source0_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [6:0] burst_adapter_001_source0_channel;                                                                   // burst_adapter_001:source0_channel -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                               // burst_adapter_002:source0_endofpacket -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                     // burst_adapter_002:source0_valid -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                             // burst_adapter_002:source0_startofpacket -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [109:0] burst_adapter_002_source0_data;                                                                      // burst_adapter_002:source0_data -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                     // wrapper_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire    [6:0] burst_adapter_002_source0_channel;                                                                   // burst_adapter_002:source0_channel -> wrapper_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                               // burst_adapter_003:source0_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                     // burst_adapter_003:source0_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                             // burst_adapter_003:source0_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [109:0] burst_adapter_003_source0_data;                                                                      // burst_adapter_003:source0_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire    [6:0] burst_adapter_003_source0_channel;                                                                   // burst_adapter_003:source0_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_004_source0_endofpacket;                                                               // burst_adapter_004:source0_endofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_004_source0_valid;                                                                     // burst_adapter_004:source0_valid -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_004_source0_startofpacket;                                                             // burst_adapter_004:source0_startofpacket -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [109:0] burst_adapter_004_source0_data;                                                                      // burst_adapter_004:source0_data -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_004_source0_ready;                                                                     // mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire    [6:0] burst_adapter_004_source0_channel;                                                                   // burst_adapter_004:source0_channel -> mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_003:reset, crosser:in_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, crosser_007:in_reset, crosser_008:out_reset, crosser_009:out_reset, crosser_010:out_reset, crosser_011:out_reset, crosser_012:out_reset, crosser_013:out_reset, dma:system_reset_n, dma_control_port_slave_translator:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_read_master_translator:reset, dma_read_master_translator_avalon_universal_master_0_agent:reset, dma_write_master_translator:reset, dma_write_master_translator_avalon_universal_master_0_agent:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_005:reset, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, limiter_002:reset, mm_clock_crossing_bridge_io:m0_reset, mm_clock_crossing_bridge_io_m0_translator:reset, mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent:reset, nios2_qsys:reset_n, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory:reset, onchip_memory_s1_translator:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ppl_mem_reader:reset, ppl_mem_reader_avalon_master_translator:reset, ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_005:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, wrapper_0:reset, wrapper_0_s0_translator:reset, wrapper_0_s0_translator_avalon_universal_slave_0_agent:reset, wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_reset_out_reset_req;                                                                  // rst_controller:reset_req -> onchip_memory:reset_req
	wire          rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> [burst_adapter_004:reset, button:reset_n, button_s1_translator:reset, button_s1_translator_avalon_universal_slave_0_agent:reset, button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:out_reset, crosser_008:in_reset, crosser_009:in_reset, crosser_010:in_reset, crosser_011:in_reset, crosser_012:in_reset, crosser_013:in_reset, ddr2_i2c_scl:reset_n, ddr2_i2c_scl_s1_translator:reset, ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ddr2_i2c_sda:reset_n, ddr2_i2c_sda_s1_translator:reset, ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, irq_synchronizer:receiver_reset, led:reset_n, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, mm_clock_crossing_bridge_io:s0_reset, mm_clock_crossing_bridge_io_s0_translator:reset, mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent:reset, mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_002_reset_out_reset;                                                                  // rst_controller_002:reset_out -> [cmd_xbar_mux_004:reset, id_router_004:reset, mem_if_ddr2_emif_avl_translator:reset, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:reset, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_004:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire          mem_if_ddr2_emif_afi_reset_reset;                                                                    // mem_if_ddr2_emif:afi_reset_n -> rst_controller_002:reset_in0
	wire          cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [109:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [6:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [109:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [6:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [109:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [6:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                                     // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                           // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                   // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [109:0] cmd_xbar_demux_src3_data;                                                                            // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire    [6:0] cmd_xbar_demux_src3_channel;                                                                         // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                           // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [109:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [6:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [109:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [6:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [109:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_003:sink1_data
	wire    [6:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [109:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> burst_adapter_003:sink0_data
	wire    [6:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> burst_adapter_003:sink0_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [109:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [6:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [109:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [6:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [109:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [6:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [109:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [6:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [109:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [6:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [109:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [6:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                 // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                       // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                               // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [109:0] rsp_xbar_demux_003_src1_data;                                                                        // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink2_data
	wire    [6:0] rsp_xbar_demux_003_src1_channel;                                                                     // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [109:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [6:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_005:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                         // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                       // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [109:0] limiter_cmd_src_data;                                                                                // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [6:0] limiter_cmd_src_channel;                                                                             // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [109:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [6:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                              // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                     // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                   // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [109:0] limiter_001_cmd_src_data;                                                                            // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire    [6:0] limiter_001_cmd_src_channel;                                                                         // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [109:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire    [6:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                          // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                     // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                           // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                   // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [91:0] addr_router_002_src_data;                                                                            // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [6:0] addr_router_002_src_channel;                                                                         // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                           // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          width_adapter_005_src_ready;                                                                         // dma_read_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_005:out_ready
	wire          addr_router_003_src_endofpacket;                                                                     // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                           // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                   // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [91:0] addr_router_003_src_data;                                                                            // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [6:0] addr_router_003_src_channel;                                                                         // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                           // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          width_adapter_006_src_ready;                                                                         // dma_write_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_006:out_ready
	wire          addr_router_004_src_endofpacket;                                                                     // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                           // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                   // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [109:0] addr_router_004_src_data;                                                                            // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire    [6:0] addr_router_004_src_channel;                                                                         // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                           // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          width_adapter_007_src_ready;                                                                         // ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_007:out_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [109:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> burst_adapter:sink0_data
	wire    [6:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_src_ready;                                                                              // burst_adapter:sink0_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [109:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [6:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [109:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> burst_adapter_001:sink0_data
	wire    [6:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                          // burst_adapter_001:sink0_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [109:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [6:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src2_ready;                                                                           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire          id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [109:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [6:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                    // cmd_xbar_mux_003:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                          // cmd_xbar_mux_003:src_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                  // cmd_xbar_mux_003:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [109:0] cmd_xbar_mux_003_src_data;                                                                           // cmd_xbar_mux_003:src_data -> burst_adapter_002:sink0_data
	wire    [6:0] cmd_xbar_mux_003_src_channel;                                                                        // cmd_xbar_mux_003:src_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                          // burst_adapter_002:sink0_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [109:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [6:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                    // cmd_xbar_mux_004:src_endofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                          // cmd_xbar_mux_004:src_valid -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                  // cmd_xbar_mux_004:src_startofpacket -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [361:0] cmd_xbar_mux_004_src_data;                                                                           // cmd_xbar_mux_004:src_data -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire    [6:0] cmd_xbar_mux_004_src_channel;                                                                        // cmd_xbar_mux_004:src_channel -> mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                          // mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [361:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [6:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                       // burst_adapter_003:sink0_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [109:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [6:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          crosser_out_ready;                                                                                   // burst_adapter_004:sink0_ready -> crosser:out_ready
	wire          id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [109:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [6:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                     // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                   // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire   [80:0] limiter_002_cmd_src_data;                                                                            // limiter_002:cmd_src_data -> cmd_xbar_demux_005:sink_data
	wire    [5:0] limiter_002_cmd_src_channel;                                                                         // limiter_002:cmd_src_channel -> cmd_xbar_demux_005:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                           // cmd_xbar_demux_005:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_005_src_endofpacket;                                                                    // rsp_xbar_mux_005:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_005_src_valid;                                                                          // rsp_xbar_mux_005:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_005_src_startofpacket;                                                                  // rsp_xbar_mux_005:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [80:0] rsp_xbar_mux_005_src_data;                                                                           // rsp_xbar_mux_005:src_data -> limiter_002:rsp_sink_data
	wire    [5:0] rsp_xbar_mux_005_src_channel;                                                                        // rsp_xbar_mux_005:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_005_src_ready;                                                                          // limiter_002:rsp_sink_ready -> rsp_xbar_mux_005:src_ready
	wire          crosser_002_out_ready;                                                                               // button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire          id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [80:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [5:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          crosser_003_out_ready;                                                                               // led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_003:out_ready
	wire          id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [80:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [5:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          crosser_004_out_ready;                                                                               // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_004:out_ready
	wire          id_router_009_src_endofpacket;                                                                       // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                             // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                     // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [80:0] id_router_009_src_data;                                                                              // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire    [5:0] id_router_009_src_channel;                                                                           // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                             // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          crosser_005_out_ready;                                                                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_005:out_ready
	wire          id_router_010_src_endofpacket;                                                                       // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                             // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                     // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [80:0] id_router_010_src_data;                                                                              // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire    [5:0] id_router_010_src_channel;                                                                           // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                             // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          crosser_006_out_ready;                                                                               // ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_006:out_ready
	wire          id_router_011_src_endofpacket;                                                                       // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                             // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                     // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [80:0] id_router_011_src_data;                                                                              // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire    [5:0] id_router_011_src_channel;                                                                           // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                             // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          crosser_007_out_ready;                                                                               // ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_007:out_ready
	wire          id_router_012_src_endofpacket;                                                                       // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                             // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                     // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [80:0] id_router_012_src_data;                                                                              // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire    [5:0] id_router_012_src_channel;                                                                           // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                             // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> width_adapter:in_startofpacket
	wire  [109:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> width_adapter:in_data
	wire    [6:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_demux_001:src3_ready
	wire          width_adapter_src_endofpacket;                                                                       // width_adapter:out_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                             // width_adapter:out_valid -> cmd_xbar_mux_004:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                     // width_adapter:out_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [361:0] width_adapter_src_data;                                                                              // width_adapter:out_data -> cmd_xbar_mux_004:sink0_data
	wire          width_adapter_src_ready;                                                                             // cmd_xbar_mux_004:sink0_ready -> width_adapter:out_ready
	wire    [6:0] width_adapter_src_channel;                                                                           // width_adapter:out_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                 // cmd_xbar_demux_002:src0_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                       // cmd_xbar_demux_002:src0_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                               // cmd_xbar_demux_002:src0_startofpacket -> width_adapter_001:in_startofpacket
	wire   [91:0] cmd_xbar_demux_002_src0_data;                                                                        // cmd_xbar_demux_002:src0_data -> width_adapter_001:in_data
	wire    [6:0] cmd_xbar_demux_002_src0_channel;                                                                     // cmd_xbar_demux_002:src0_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                       // width_adapter_001:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          width_adapter_001_src_endofpacket;                                                                   // width_adapter_001:out_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          width_adapter_001_src_valid;                                                                         // width_adapter_001:out_valid -> cmd_xbar_mux_004:sink1_valid
	wire          width_adapter_001_src_startofpacket;                                                                 // width_adapter_001:out_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [361:0] width_adapter_001_src_data;                                                                          // width_adapter_001:out_data -> cmd_xbar_mux_004:sink1_data
	wire          width_adapter_001_src_ready;                                                                         // cmd_xbar_mux_004:sink1_ready -> width_adapter_001:out_ready
	wire    [6:0] width_adapter_001_src_channel;                                                                       // width_adapter_001:out_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                 // cmd_xbar_demux_003:src0_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                       // cmd_xbar_demux_003:src0_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                               // cmd_xbar_demux_003:src0_startofpacket -> width_adapter_002:in_startofpacket
	wire   [91:0] cmd_xbar_demux_003_src0_data;                                                                        // cmd_xbar_demux_003:src0_data -> width_adapter_002:in_data
	wire    [6:0] cmd_xbar_demux_003_src0_channel;                                                                     // cmd_xbar_demux_003:src0_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                       // width_adapter_002:in_ready -> cmd_xbar_demux_003:src0_ready
	wire          width_adapter_002_src_endofpacket;                                                                   // width_adapter_002:out_endofpacket -> cmd_xbar_mux_004:sink2_endofpacket
	wire          width_adapter_002_src_valid;                                                                         // width_adapter_002:out_valid -> cmd_xbar_mux_004:sink2_valid
	wire          width_adapter_002_src_startofpacket;                                                                 // width_adapter_002:out_startofpacket -> cmd_xbar_mux_004:sink2_startofpacket
	wire  [361:0] width_adapter_002_src_data;                                                                          // width_adapter_002:out_data -> cmd_xbar_mux_004:sink2_data
	wire          width_adapter_002_src_ready;                                                                         // cmd_xbar_mux_004:sink2_ready -> width_adapter_002:out_ready
	wire    [6:0] width_adapter_002_src_channel;                                                                       // width_adapter_002:out_channel -> cmd_xbar_mux_004:sink2_channel
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                 // cmd_xbar_demux_004:src0_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                       // cmd_xbar_demux_004:src0_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                               // cmd_xbar_demux_004:src0_startofpacket -> width_adapter_003:in_startofpacket
	wire  [109:0] cmd_xbar_demux_004_src0_data;                                                                        // cmd_xbar_demux_004:src0_data -> width_adapter_003:in_data
	wire    [6:0] cmd_xbar_demux_004_src0_channel;                                                                     // cmd_xbar_demux_004:src0_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                       // width_adapter_003:in_ready -> cmd_xbar_demux_004:src0_ready
	wire          width_adapter_003_src_endofpacket;                                                                   // width_adapter_003:out_endofpacket -> cmd_xbar_mux_004:sink3_endofpacket
	wire          width_adapter_003_src_valid;                                                                         // width_adapter_003:out_valid -> cmd_xbar_mux_004:sink3_valid
	wire          width_adapter_003_src_startofpacket;                                                                 // width_adapter_003:out_startofpacket -> cmd_xbar_mux_004:sink3_startofpacket
	wire  [361:0] width_adapter_003_src_data;                                                                          // width_adapter_003:out_data -> cmd_xbar_mux_004:sink3_data
	wire          width_adapter_003_src_ready;                                                                         // cmd_xbar_mux_004:sink3_ready -> width_adapter_003:out_ready
	wire    [6:0] width_adapter_003_src_channel;                                                                       // width_adapter_003:out_channel -> cmd_xbar_mux_004:sink3_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> width_adapter_004:in_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> width_adapter_004:in_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> width_adapter_004:in_startofpacket
	wire  [361:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> width_adapter_004:in_data
	wire    [6:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> width_adapter_004:in_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                       // width_adapter_004:in_ready -> rsp_xbar_demux_004:src0_ready
	wire          width_adapter_004_src_endofpacket;                                                                   // width_adapter_004:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          width_adapter_004_src_valid;                                                                         // width_adapter_004:out_valid -> rsp_xbar_mux_001:sink3_valid
	wire          width_adapter_004_src_startofpacket;                                                                 // width_adapter_004:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [109:0] width_adapter_004_src_data;                                                                          // width_adapter_004:out_data -> rsp_xbar_mux_001:sink3_data
	wire          width_adapter_004_src_ready;                                                                         // rsp_xbar_mux_001:sink3_ready -> width_adapter_004:out_ready
	wire    [6:0] width_adapter_004_src_channel;                                                                       // width_adapter_004:out_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                 // rsp_xbar_demux_004:src1_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                       // rsp_xbar_demux_004:src1_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                               // rsp_xbar_demux_004:src1_startofpacket -> width_adapter_005:in_startofpacket
	wire  [361:0] rsp_xbar_demux_004_src1_data;                                                                        // rsp_xbar_demux_004:src1_data -> width_adapter_005:in_data
	wire    [6:0] rsp_xbar_demux_004_src1_channel;                                                                     // rsp_xbar_demux_004:src1_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                       // width_adapter_005:in_ready -> rsp_xbar_demux_004:src1_ready
	wire          width_adapter_005_src_endofpacket;                                                                   // width_adapter_005:out_endofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_005_src_valid;                                                                         // width_adapter_005:out_valid -> dma_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_005_src_startofpacket;                                                                 // width_adapter_005:out_startofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [91:0] width_adapter_005_src_data;                                                                          // width_adapter_005:out_data -> dma_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [6:0] width_adapter_005_src_channel;                                                                       // width_adapter_005:out_channel -> dma_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src2_endofpacket;                                                                 // rsp_xbar_demux_004:src2_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_004_src2_valid;                                                                       // rsp_xbar_demux_004:src2_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_004_src2_startofpacket;                                                               // rsp_xbar_demux_004:src2_startofpacket -> width_adapter_006:in_startofpacket
	wire  [361:0] rsp_xbar_demux_004_src2_data;                                                                        // rsp_xbar_demux_004:src2_data -> width_adapter_006:in_data
	wire    [6:0] rsp_xbar_demux_004_src2_channel;                                                                     // rsp_xbar_demux_004:src2_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_004_src2_ready;                                                                       // width_adapter_006:in_ready -> rsp_xbar_demux_004:src2_ready
	wire          width_adapter_006_src_endofpacket;                                                                   // width_adapter_006:out_endofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_006_src_valid;                                                                         // width_adapter_006:out_valid -> dma_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_006_src_startofpacket;                                                                 // width_adapter_006:out_startofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [91:0] width_adapter_006_src_data;                                                                          // width_adapter_006:out_data -> dma_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [6:0] width_adapter_006_src_channel;                                                                       // width_adapter_006:out_channel -> dma_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src3_endofpacket;                                                                 // rsp_xbar_demux_004:src3_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_004_src3_valid;                                                                       // rsp_xbar_demux_004:src3_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_004_src3_startofpacket;                                                               // rsp_xbar_demux_004:src3_startofpacket -> width_adapter_007:in_startofpacket
	wire  [361:0] rsp_xbar_demux_004_src3_data;                                                                        // rsp_xbar_demux_004:src3_data -> width_adapter_007:in_data
	wire    [6:0] rsp_xbar_demux_004_src3_channel;                                                                     // rsp_xbar_demux_004:src3_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_004_src3_ready;                                                                       // width_adapter_007:in_ready -> rsp_xbar_demux_004:src3_ready
	wire          width_adapter_007_src_endofpacket;                                                                   // width_adapter_007:out_endofpacket -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_007_src_valid;                                                                         // width_adapter_007:out_valid -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_007_src_startofpacket;                                                                 // width_adapter_007:out_startofpacket -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [109:0] width_adapter_007_src_data;                                                                          // width_adapter_007:out_data -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [6:0] width_adapter_007_src_channel;                                                                       // width_adapter_007:out_channel -> ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          crosser_out_endofpacket;                                                                             // crosser:out_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire          crosser_out_valid;                                                                                   // crosser:out_valid -> burst_adapter_004:sink0_valid
	wire          crosser_out_startofpacket;                                                                           // crosser:out_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire  [109:0] crosser_out_data;                                                                                    // crosser:out_data -> burst_adapter_004:sink0_data
	wire    [6:0] crosser_out_channel;                                                                                 // crosser:out_channel -> burst_adapter_004:sink0_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> crosser:in_startofpacket
	wire  [109:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> crosser:in_data
	wire    [6:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                       // crosser:in_ready -> cmd_xbar_demux_001:src5_ready
	wire          crosser_001_out_endofpacket;                                                                         // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          crosser_001_out_valid;                                                                               // crosser_001:out_valid -> rsp_xbar_mux_001:sink5_valid
	wire          crosser_001_out_startofpacket;                                                                       // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [109:0] crosser_001_out_data;                                                                                // crosser_001:out_data -> rsp_xbar_mux_001:sink5_data
	wire    [6:0] crosser_001_out_channel;                                                                             // crosser_001:out_channel -> rsp_xbar_mux_001:sink5_channel
	wire          crosser_001_out_ready;                                                                               // rsp_xbar_mux_001:sink5_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [109:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> crosser_001:in_data
	wire    [6:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                       // crosser_001:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          crosser_002_out_endofpacket;                                                                         // crosser_002:out_endofpacket -> button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_002_out_valid;                                                                               // crosser_002:out_valid -> button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_002_out_startofpacket;                                                                       // crosser_002:out_startofpacket -> button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] crosser_002_out_data;                                                                                // crosser_002:out_data -> button_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_002_out_channel;                                                                             // crosser_002:out_channel -> button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                 // cmd_xbar_demux_005:src0_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                       // cmd_xbar_demux_005:src0_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                               // cmd_xbar_demux_005:src0_startofpacket -> crosser_002:in_startofpacket
	wire   [80:0] cmd_xbar_demux_005_src0_data;                                                                        // cmd_xbar_demux_005:src0_data -> crosser_002:in_data
	wire    [5:0] cmd_xbar_demux_005_src0_channel;                                                                     // cmd_xbar_demux_005:src0_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                       // crosser_002:in_ready -> cmd_xbar_demux_005:src0_ready
	wire          crosser_003_out_endofpacket;                                                                         // crosser_003:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_003_out_valid;                                                                               // crosser_003:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_003_out_startofpacket;                                                                       // crosser_003:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] crosser_003_out_data;                                                                                // crosser_003:out_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_003_out_channel;                                                                             // crosser_003:out_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src1_endofpacket;                                                                 // cmd_xbar_demux_005:src1_endofpacket -> crosser_003:in_endofpacket
	wire          cmd_xbar_demux_005_src1_valid;                                                                       // cmd_xbar_demux_005:src1_valid -> crosser_003:in_valid
	wire          cmd_xbar_demux_005_src1_startofpacket;                                                               // cmd_xbar_demux_005:src1_startofpacket -> crosser_003:in_startofpacket
	wire   [80:0] cmd_xbar_demux_005_src1_data;                                                                        // cmd_xbar_demux_005:src1_data -> crosser_003:in_data
	wire    [5:0] cmd_xbar_demux_005_src1_channel;                                                                     // cmd_xbar_demux_005:src1_channel -> crosser_003:in_channel
	wire          cmd_xbar_demux_005_src1_ready;                                                                       // crosser_003:in_ready -> cmd_xbar_demux_005:src1_ready
	wire          crosser_004_out_endofpacket;                                                                         // crosser_004:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_004_out_valid;                                                                               // crosser_004:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_004_out_startofpacket;                                                                       // crosser_004:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] crosser_004_out_data;                                                                                // crosser_004:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_004_out_channel;                                                                             // crosser_004:out_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src2_endofpacket;                                                                 // cmd_xbar_demux_005:src2_endofpacket -> crosser_004:in_endofpacket
	wire          cmd_xbar_demux_005_src2_valid;                                                                       // cmd_xbar_demux_005:src2_valid -> crosser_004:in_valid
	wire          cmd_xbar_demux_005_src2_startofpacket;                                                               // cmd_xbar_demux_005:src2_startofpacket -> crosser_004:in_startofpacket
	wire   [80:0] cmd_xbar_demux_005_src2_data;                                                                        // cmd_xbar_demux_005:src2_data -> crosser_004:in_data
	wire    [5:0] cmd_xbar_demux_005_src2_channel;                                                                     // cmd_xbar_demux_005:src2_channel -> crosser_004:in_channel
	wire          cmd_xbar_demux_005_src2_ready;                                                                       // crosser_004:in_ready -> cmd_xbar_demux_005:src2_ready
	wire          crosser_005_out_endofpacket;                                                                         // crosser_005:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_005_out_valid;                                                                               // crosser_005:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_005_out_startofpacket;                                                                       // crosser_005:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] crosser_005_out_data;                                                                                // crosser_005:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_005_out_channel;                                                                             // crosser_005:out_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src3_endofpacket;                                                                 // cmd_xbar_demux_005:src3_endofpacket -> crosser_005:in_endofpacket
	wire          cmd_xbar_demux_005_src3_valid;                                                                       // cmd_xbar_demux_005:src3_valid -> crosser_005:in_valid
	wire          cmd_xbar_demux_005_src3_startofpacket;                                                               // cmd_xbar_demux_005:src3_startofpacket -> crosser_005:in_startofpacket
	wire   [80:0] cmd_xbar_demux_005_src3_data;                                                                        // cmd_xbar_demux_005:src3_data -> crosser_005:in_data
	wire    [5:0] cmd_xbar_demux_005_src3_channel;                                                                     // cmd_xbar_demux_005:src3_channel -> crosser_005:in_channel
	wire          cmd_xbar_demux_005_src3_ready;                                                                       // crosser_005:in_ready -> cmd_xbar_demux_005:src3_ready
	wire          crosser_006_out_endofpacket;                                                                         // crosser_006:out_endofpacket -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_006_out_valid;                                                                               // crosser_006:out_valid -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_006_out_startofpacket;                                                                       // crosser_006:out_startofpacket -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] crosser_006_out_data;                                                                                // crosser_006:out_data -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_006_out_channel;                                                                             // crosser_006:out_channel -> ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src4_endofpacket;                                                                 // cmd_xbar_demux_005:src4_endofpacket -> crosser_006:in_endofpacket
	wire          cmd_xbar_demux_005_src4_valid;                                                                       // cmd_xbar_demux_005:src4_valid -> crosser_006:in_valid
	wire          cmd_xbar_demux_005_src4_startofpacket;                                                               // cmd_xbar_demux_005:src4_startofpacket -> crosser_006:in_startofpacket
	wire   [80:0] cmd_xbar_demux_005_src4_data;                                                                        // cmd_xbar_demux_005:src4_data -> crosser_006:in_data
	wire    [5:0] cmd_xbar_demux_005_src4_channel;                                                                     // cmd_xbar_demux_005:src4_channel -> crosser_006:in_channel
	wire          cmd_xbar_demux_005_src4_ready;                                                                       // crosser_006:in_ready -> cmd_xbar_demux_005:src4_ready
	wire          crosser_007_out_endofpacket;                                                                         // crosser_007:out_endofpacket -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_007_out_valid;                                                                               // crosser_007:out_valid -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_007_out_startofpacket;                                                                       // crosser_007:out_startofpacket -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [80:0] crosser_007_out_data;                                                                                // crosser_007:out_data -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] crosser_007_out_channel;                                                                             // crosser_007:out_channel -> ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src5_endofpacket;                                                                 // cmd_xbar_demux_005:src5_endofpacket -> crosser_007:in_endofpacket
	wire          cmd_xbar_demux_005_src5_valid;                                                                       // cmd_xbar_demux_005:src5_valid -> crosser_007:in_valid
	wire          cmd_xbar_demux_005_src5_startofpacket;                                                               // cmd_xbar_demux_005:src5_startofpacket -> crosser_007:in_startofpacket
	wire   [80:0] cmd_xbar_demux_005_src5_data;                                                                        // cmd_xbar_demux_005:src5_data -> crosser_007:in_data
	wire    [5:0] cmd_xbar_demux_005_src5_channel;                                                                     // cmd_xbar_demux_005:src5_channel -> crosser_007:in_channel
	wire          cmd_xbar_demux_005_src5_ready;                                                                       // crosser_007:in_ready -> cmd_xbar_demux_005:src5_ready
	wire          crosser_008_out_endofpacket;                                                                         // crosser_008:out_endofpacket -> rsp_xbar_mux_005:sink0_endofpacket
	wire          crosser_008_out_valid;                                                                               // crosser_008:out_valid -> rsp_xbar_mux_005:sink0_valid
	wire          crosser_008_out_startofpacket;                                                                       // crosser_008:out_startofpacket -> rsp_xbar_mux_005:sink0_startofpacket
	wire   [80:0] crosser_008_out_data;                                                                                // crosser_008:out_data -> rsp_xbar_mux_005:sink0_data
	wire    [5:0] crosser_008_out_channel;                                                                             // crosser_008:out_channel -> rsp_xbar_mux_005:sink0_channel
	wire          crosser_008_out_ready;                                                                               // rsp_xbar_mux_005:sink0_ready -> crosser_008:out_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> crosser_008:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> crosser_008:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> crosser_008:in_startofpacket
	wire   [80:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> crosser_008:in_data
	wire    [5:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> crosser_008:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                       // crosser_008:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          crosser_009_out_endofpacket;                                                                         // crosser_009:out_endofpacket -> rsp_xbar_mux_005:sink1_endofpacket
	wire          crosser_009_out_valid;                                                                               // crosser_009:out_valid -> rsp_xbar_mux_005:sink1_valid
	wire          crosser_009_out_startofpacket;                                                                       // crosser_009:out_startofpacket -> rsp_xbar_mux_005:sink1_startofpacket
	wire   [80:0] crosser_009_out_data;                                                                                // crosser_009:out_data -> rsp_xbar_mux_005:sink1_data
	wire    [5:0] crosser_009_out_channel;                                                                             // crosser_009:out_channel -> rsp_xbar_mux_005:sink1_channel
	wire          crosser_009_out_ready;                                                                               // rsp_xbar_mux_005:sink1_ready -> crosser_009:out_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> crosser_009:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> crosser_009:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> crosser_009:in_startofpacket
	wire   [80:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> crosser_009:in_data
	wire    [5:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> crosser_009:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                       // crosser_009:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          crosser_010_out_endofpacket;                                                                         // crosser_010:out_endofpacket -> rsp_xbar_mux_005:sink2_endofpacket
	wire          crosser_010_out_valid;                                                                               // crosser_010:out_valid -> rsp_xbar_mux_005:sink2_valid
	wire          crosser_010_out_startofpacket;                                                                       // crosser_010:out_startofpacket -> rsp_xbar_mux_005:sink2_startofpacket
	wire   [80:0] crosser_010_out_data;                                                                                // crosser_010:out_data -> rsp_xbar_mux_005:sink2_data
	wire    [5:0] crosser_010_out_channel;                                                                             // crosser_010:out_channel -> rsp_xbar_mux_005:sink2_channel
	wire          crosser_010_out_ready;                                                                               // rsp_xbar_mux_005:sink2_ready -> crosser_010:out_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                 // rsp_xbar_demux_009:src0_endofpacket -> crosser_010:in_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                       // rsp_xbar_demux_009:src0_valid -> crosser_010:in_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                               // rsp_xbar_demux_009:src0_startofpacket -> crosser_010:in_startofpacket
	wire   [80:0] rsp_xbar_demux_009_src0_data;                                                                        // rsp_xbar_demux_009:src0_data -> crosser_010:in_data
	wire    [5:0] rsp_xbar_demux_009_src0_channel;                                                                     // rsp_xbar_demux_009:src0_channel -> crosser_010:in_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                       // crosser_010:in_ready -> rsp_xbar_demux_009:src0_ready
	wire          crosser_011_out_endofpacket;                                                                         // crosser_011:out_endofpacket -> rsp_xbar_mux_005:sink3_endofpacket
	wire          crosser_011_out_valid;                                                                               // crosser_011:out_valid -> rsp_xbar_mux_005:sink3_valid
	wire          crosser_011_out_startofpacket;                                                                       // crosser_011:out_startofpacket -> rsp_xbar_mux_005:sink3_startofpacket
	wire   [80:0] crosser_011_out_data;                                                                                // crosser_011:out_data -> rsp_xbar_mux_005:sink3_data
	wire    [5:0] crosser_011_out_channel;                                                                             // crosser_011:out_channel -> rsp_xbar_mux_005:sink3_channel
	wire          crosser_011_out_ready;                                                                               // rsp_xbar_mux_005:sink3_ready -> crosser_011:out_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                 // rsp_xbar_demux_010:src0_endofpacket -> crosser_011:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                       // rsp_xbar_demux_010:src0_valid -> crosser_011:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                               // rsp_xbar_demux_010:src0_startofpacket -> crosser_011:in_startofpacket
	wire   [80:0] rsp_xbar_demux_010_src0_data;                                                                        // rsp_xbar_demux_010:src0_data -> crosser_011:in_data
	wire    [5:0] rsp_xbar_demux_010_src0_channel;                                                                     // rsp_xbar_demux_010:src0_channel -> crosser_011:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                       // crosser_011:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          crosser_012_out_endofpacket;                                                                         // crosser_012:out_endofpacket -> rsp_xbar_mux_005:sink4_endofpacket
	wire          crosser_012_out_valid;                                                                               // crosser_012:out_valid -> rsp_xbar_mux_005:sink4_valid
	wire          crosser_012_out_startofpacket;                                                                       // crosser_012:out_startofpacket -> rsp_xbar_mux_005:sink4_startofpacket
	wire   [80:0] crosser_012_out_data;                                                                                // crosser_012:out_data -> rsp_xbar_mux_005:sink4_data
	wire    [5:0] crosser_012_out_channel;                                                                             // crosser_012:out_channel -> rsp_xbar_mux_005:sink4_channel
	wire          crosser_012_out_ready;                                                                               // rsp_xbar_mux_005:sink4_ready -> crosser_012:out_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                 // rsp_xbar_demux_011:src0_endofpacket -> crosser_012:in_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                       // rsp_xbar_demux_011:src0_valid -> crosser_012:in_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                               // rsp_xbar_demux_011:src0_startofpacket -> crosser_012:in_startofpacket
	wire   [80:0] rsp_xbar_demux_011_src0_data;                                                                        // rsp_xbar_demux_011:src0_data -> crosser_012:in_data
	wire    [5:0] rsp_xbar_demux_011_src0_channel;                                                                     // rsp_xbar_demux_011:src0_channel -> crosser_012:in_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                       // crosser_012:in_ready -> rsp_xbar_demux_011:src0_ready
	wire          crosser_013_out_endofpacket;                                                                         // crosser_013:out_endofpacket -> rsp_xbar_mux_005:sink5_endofpacket
	wire          crosser_013_out_valid;                                                                               // crosser_013:out_valid -> rsp_xbar_mux_005:sink5_valid
	wire          crosser_013_out_startofpacket;                                                                       // crosser_013:out_startofpacket -> rsp_xbar_mux_005:sink5_startofpacket
	wire   [80:0] crosser_013_out_data;                                                                                // crosser_013:out_data -> rsp_xbar_mux_005:sink5_data
	wire    [5:0] crosser_013_out_channel;                                                                             // crosser_013:out_channel -> rsp_xbar_mux_005:sink5_channel
	wire          crosser_013_out_ready;                                                                               // rsp_xbar_mux_005:sink5_ready -> crosser_013:out_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                 // rsp_xbar_demux_012:src0_endofpacket -> crosser_013:in_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                       // rsp_xbar_demux_012:src0_valid -> crosser_013:in_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                               // rsp_xbar_demux_012:src0_startofpacket -> crosser_013:in_startofpacket
	wire   [80:0] rsp_xbar_demux_012_src0_data;                                                                        // rsp_xbar_demux_012:src0_data -> crosser_013:in_data
	wire    [5:0] rsp_xbar_demux_012_src0_channel;                                                                     // rsp_xbar_demux_012:src0_channel -> crosser_013:in_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                       // crosser_013:in_ready -> rsp_xbar_demux_012:src0_ready
	wire    [6:0] limiter_cmd_valid_data;                                                                              // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [6:0] limiter_001_cmd_valid_data;                                                                          // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire    [5:0] limiter_002_cmd_valid_data;                                                                          // limiter_002:cmd_src_valid -> cmd_xbar_demux_005:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                            // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver2_irq;                                                                            // dma:dma_ctl_irq -> irq_mapper:receiver2_irq
	wire   [31:0] nios2_qsys_d_irq_irq;                                                                                // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire          irq_mapper_receiver1_irq;                                                                            // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                       // timer:irq -> irq_synchronizer:receiver_irq

	DE4_QSYS_onchip_memory onchip_memory (
		.clk        (mem_if_ddr2_emif_afi_clk_clk),                               //   clk1.clk
		.address    (onchip_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                          //       .reset_req
	);

	DE4_QSYS_mem_if_ddr2_emif mem_if_ddr2_emif (
		.pll_ref_clk        (clk_clk),                                                                //      pll_ref_clk.clk
		.global_reset_n     (reset_reset_n),                                                          //     global_reset.reset_n
		.soft_reset_n       (reset_reset_n),                                                          //       soft_reset.reset_n
		.afi_clk            (mem_if_ddr2_emif_afi_clk_clk),                                           //          afi_clk.clk
		.afi_half_clk       (),                                                                       //     afi_half_clk.clk
		.afi_reset_n        (mem_if_ddr2_emif_afi_reset_reset),                                       //        afi_reset.reset_n
		.afi_reset_export_n (),                                                                       // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                                           //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                                          //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                                          //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                                        //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                                         //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                                        //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                                          //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                                       //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                                       //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                                        //                 .mem_we_n
		.mem_dq             (memory_mem_dq),                                                          //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                                         //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                                       //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                                         //                 .mem_odt
		.avl_ready          (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_address),            //                 .address
		.avl_rdata_valid    (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdata),           //                 .readdata
		.avl_wdata          (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_writedata),          //                 .writedata
		.avl_be             (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_byteenable),         //                 .byteenable
		.avl_read_req       (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_read),               //                 .read
		.avl_write_req      (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_write),              //                 .write
		.avl_size           (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_burstcount),         //                 .burstcount
		.local_init_done    (mem_if_ddr2_emif_status_local_init_done),                                //           status.local_init_done
		.local_cal_success  (mem_if_ddr2_emif_status_local_cal_success),                              //                 .local_cal_success
		.local_cal_fail     (mem_if_ddr2_emif_status_local_cal_fail),                                 //                 .local_cal_fail
		.oct_rdn            (oct_rdn),                                                                //              oct.rdn
		.oct_rup            (oct_rup)                                                                 //                 .rup
	);

	DE4_QSYS_nios2_qsys nios2_qsys (
		.clk                                   (mem_if_ddr2_emif_afi_clk_clk),                                            //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                         //                   reset_n.reset_n
		.d_address                             (nios2_qsys_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                                        //                          .writedata
		.d_burstcount                          (nios2_qsys_data_master_burstcount),                                       //                          .burstcount
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                                        //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                         // custom_instruction_master.readra
	);

	DE4_QSYS_jtag_uart jtag_uart (
		.clk            (mem_if_ddr2_emif_afi_clk_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	DE4_QSYS_sysid sysid (
		.clock    (clk_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	DE4_QSYS_timer timer (
		.clk        (clk_clk),                                            //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                       //   irq.irq
	);

	DE4_QSYS_led led (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                        // external_connection.export
	);

	DE4_QSYS_button button (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address  (button_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (button_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (button_export)                                      // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_io (
		.m0_clk           (mem_if_ddr2_emif_afi_clk_clk),                                                //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                                              // m0_reset.reset
		.s0_clk           (clk_clk),                                                                     //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                          // s0_reset.reset
		.s0_waitrequest   (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_io_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_io_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_io_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_io_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_io_m0_writedata),                                    //         .writedata
		.m0_address       (mm_clock_crossing_bridge_io_m0_address),                                      //         .address
		.m0_write         (mm_clock_crossing_bridge_io_m0_write),                                        //         .write
		.m0_read          (mm_clock_crossing_bridge_io_m0_read),                                         //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_io_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_io_m0_debugaccess)                                   //         .debugaccess
	);

	DE4_QSYS_ddr2_i2c_scl ddr2_i2c_scl (
		.clk        (clk_clk),                                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address    (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ddr2_i2c_scl_export)                                        // external_connection.export
	);

	DE4_QSYS_ddr2_i2c_sda ddr2_i2c_sda (
		.clk        (clk_clk),                                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                       //               reset.reset_n
		.address    (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (ddr2_i2c_sda_export)                                        // external_connection.export
	);

	DE4_QSYS_dma dma (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                     //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                  //              reset.reset_n
		.dma_ctl_address    (dma_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver2_irq),                                         //                irq.irq
		.read_address       (dma_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_read_master_waitrequest),                                      //                   .waitrequest
		.read_burstcount    (dma_read_master_burstcount),                                       //                   .burstcount
		.write_address      (dma_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_write_master_byteenable),                                      //                   .byteenable
		.write_burstcount   (dma_write_master_burstcount)                                       //                   .burstcount
	);

	latency_aware_read_master #(
		.DATAWIDTH       (32),
		.BYTEENABLEWIDTH (4),
		.ADDRESSWIDTH    (32),
		.FIFODEPTH       (32),
		.FIFODEPTH_LOG2  (5),
		.FIFOUSEMEMORY   (1)
	) ppl_mem_reader (
		.clk                        (mem_if_ddr2_emif_afi_clk_clk),               //         clock.clk
		.reset                      (rst_controller_reset_out_reset),             //         reset.reset
		.master_address             (ppl_mem_reader_avalon_master_address),       // avalon_master.address
		.master_read                (ppl_mem_reader_avalon_master_read),          //              .read
		.master_byteenable          (ppl_mem_reader_avalon_master_byteenable),    //              .byteenable
		.master_readdata            (ppl_mem_reader_avalon_master_readdata),      //              .readdata
		.master_readdatavalid       (ppl_mem_reader_avalon_master_readdatavalid), //              .readdatavalid
		.master_waitrequest         (ppl_mem_reader_avalon_master_waitrequest),   //              .waitrequest
		.coe_control_fixed_location (wrapper_0_control_fixed_location),           //       control.export
		.coe_control_read_base      (wrapper_0_control_read_base),                //              .export
		.coe_control_read_length    (wrapper_0_control_read_length),              //              .export
		.coe_control_go             (wrapper_0_control_go),                       //              .export
		.coe_control_done           (ppl_mem_reader_control_done),                //              .export
		.coe_control_early_done     (ppl_mem_reader_control_early_done),          //              .export
		.coe_user_read_buffer       (wrapper_0_user_read_buffer),                 //          user.export
		.coe_user_data_available    (ppl_mem_reader_user_data_available),         //              .export
		.coe_user_buffer_data       (ppl_mem_reader_user_buffer_data)             //              .export
	);

	rbm_demo #(
		.DATAWIDTH     (32),
		.ADDRESS_WIDTH (32)
	) wrapper_0 (
		.clk                        (mem_if_ddr2_emif_afi_clk_clk),                              //   clock.clk
		.reset                      (rst_controller_reset_out_reset),                            //   reset.reset
		.avs_s0_address             (wrapper_0_s0_translator_avalon_anti_slave_0_address),       //      s0.address
		.avs_s0_read                (wrapper_0_s0_translator_avalon_anti_slave_0_read),          //        .read
		.avs_s0_write               (wrapper_0_s0_translator_avalon_anti_slave_0_write),         //        .write
		.avs_s0_readdata            (wrapper_0_s0_translator_avalon_anti_slave_0_readdata),      //        .readdata
		.avs_s0_readdatavalid       (wrapper_0_s0_translator_avalon_anti_slave_0_readdatavalid), //        .readdatavalid
		.avs_s0_writedata           (wrapper_0_s0_translator_avalon_anti_slave_0_writedata),     //        .writedata
		.coe_user_data_available    (ppl_mem_reader_user_data_available),                        //    user.export
		.coe_user_read_buffer       (wrapper_0_user_read_buffer),                                //        .export
		.coe_user_buffer_data       (ppl_mem_reader_user_buffer_data),                           //        .export
		.coe_control_fixed_location (wrapper_0_control_fixed_location),                          // control.export
		.coe_control_read_base      (wrapper_0_control_read_base),                               //        .export
		.coe_control_read_length    (wrapper_0_control_read_length),                             //        .export
		.coe_control_go             (wrapper_0_control_go),                                      //        .export
		.coe_control_done           (ppl_mem_reader_control_done),                               //        .export
		.coe_control_early_done     (ppl_mem_reader_control_early_done)                          //        .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (31),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_instruction_master_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                             //               (terminated)
		.av_byteenable            (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                                             //               (terminated)
		.av_write                 (1'b0),                                                                             //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock                  (1'b0),                                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                                             //               (terminated)
		.uav_clken                (),                                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                                             //               (terminated)
		.uav_response             (2'b00),                                                                            //               (terminated)
		.av_response              (),                                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (31),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (6),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_data_master_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                              //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (nios2_qsys_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (nios2_qsys_data_master_burstcount),                                         //                          .burstcount
		.av_byteenable            (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_qsys_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_read_master_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address              (dma_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_read_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dma_read_master_burstcount),                                         //                          .burstcount
		.av_chipselect            (dma_read_master_chipselect),                                         //                          .chipselect
		.av_read                  (~dma_read_master_read),                                              //                          .read
		.av_readdata              (dma_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (dma_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable            (2'b11),                                                              //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_write                 (1'b0),                                                               //               (terminated)
		.av_writedata             (16'b0000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_write_master_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                        //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address              (dma_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_write_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dma_write_master_burstcount),                                         //                          .burstcount
		.av_byteenable            (dma_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect            (dma_write_master_chipselect),                                         //                          .chipselect
		.av_write                 (~dma_write_master_write),                                             //                          .write
		.av_writedata             (dma_write_master_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                                //               (terminated)
		.av_begintransfer         (1'b0),                                                                //               (terminated)
		.av_read                  (1'b0),                                                                //               (terminated)
		.av_readdata              (),                                                                    //               (terminated)
		.av_readdatavalid         (),                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                //               (terminated)
		.av_debugaccess           (1'b0),                                                                //               (terminated)
		.uav_clken                (),                                                                    //               (terminated)
		.av_clken                 (1'b1),                                                                //               (terminated)
		.uav_response             (2'b00),                                                               //               (terminated)
		.av_response              (),                                                                    //               (terminated)
		.uav_writeresponserequest (),                                                                    //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                //               (terminated)
		.av_writeresponsevalid    ()                                                                     //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ppl_mem_reader_avalon_master_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                    //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                  //                     reset.reset
		.uav_address              (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (ppl_mem_reader_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (ppl_mem_reader_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (ppl_mem_reader_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (ppl_mem_reader_avalon_master_read),                                               //                          .read
		.av_readdata              (ppl_mem_reader_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (ppl_mem_reader_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                            //               (terminated)
		.av_begintransfer         (1'b0),                                                                            //               (terminated)
		.av_chipselect            (1'b0),                                                                            //               (terminated)
		.av_write                 (1'b0),                                                                            //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                            //               (terminated)
		.av_lock                  (1'b0),                                                                            //               (terminated)
		.av_debugaccess           (1'b0),                                                                            //               (terminated)
		.uav_clken                (),                                                                                //               (terminated)
		.av_clken                 (1'b1),                                                                            //               (terminated)
		.uav_response             (2'b00),                                                                           //               (terminated)
		.av_response              (),                                                                                //               (terminated)
		.uav_writeresponserequest (),                                                                                //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                            //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                            //               (terminated)
		.av_writeresponsevalid    ()                                                                                 //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_jtag_debug_module_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_chipselect            (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s1_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (31),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_control_port_slave_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dma_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dma_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                  //              (terminated)
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) wrapper_0_s0_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (wrapper_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (wrapper_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (wrapper_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (wrapper_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (wrapper_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_readdatavalid         (wrapper_0_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_chipselect            (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (256),
		.UAV_DATA_W                     (256),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (32),
		.UAV_BYTEENABLE_W               (32),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (8),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (32),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mem_if_ddr2_emif_avl_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                              //                    reset.reset
		.uav_address              (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~mem_if_ddr2_emif_avl_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_chipselect            (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mm_clock_crossing_bridge_io_s0_translator (
		.clk                      (clk_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (mm_clock_crossing_bridge_io_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) mm_clock_crossing_bridge_io_m0_translator (
		.clk                      (mem_if_ddr2_emif_afi_clk_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                     reset.reset
		.uav_address              (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (mm_clock_crossing_bridge_io_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (mm_clock_crossing_bridge_io_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (mm_clock_crossing_bridge_io_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (mm_clock_crossing_bridge_io_m0_byteenable),                                         //                          .byteenable
		.av_read                  (mm_clock_crossing_bridge_io_m0_read),                                               //                          .read
		.av_readdata              (mm_clock_crossing_bridge_io_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (mm_clock_crossing_bridge_io_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (mm_clock_crossing_bridge_io_m0_write),                                              //                          .write
		.av_writedata             (mm_clock_crossing_bridge_io_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (mm_clock_crossing_bridge_io_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                              //               (terminated)
		.av_begintransfer         (1'b0),                                                                              //               (terminated)
		.av_chipselect            (1'b0),                                                                              //               (terminated)
		.av_lock                  (1'b0),                                                                              //               (terminated)
		.uav_clken                (),                                                                                  //               (terminated)
		.av_clken                 (1'b1),                                                                              //               (terminated)
		.uav_response             (2'b00),                                                                             //               (terminated)
		.av_response              (),                                                                                  //               (terminated)
		.uav_writeresponserequest (),                                                                                  //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                              //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                              //               (terminated)
		.av_writeresponsevalid    ()                                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (button_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (button_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                     //              (terminated)
		.av_read                  (),                                                                     //              (terminated)
		.av_writedata             (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_chipselect            (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_i2c_scl_s1_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ddr2_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_i2c_sda_s1_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ddr2_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_BEGIN_BURST           (92),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_THREAD_ID_H           (100),
		.PKT_THREAD_ID_L           (100),
		.PKT_CACHE_H               (107),
		.PKT_CACHE_L               (104),
		.PKT_DATA_SIDEBAND_H       (91),
		.PKT_DATA_SIDEBAND_L       (91),
		.PKT_QOS_H                 (93),
		.PKT_QOS_L                 (93),
		.PKT_ADDR_SIDEBAND_H       (90),
		.PKT_ADDR_SIDEBAND_L       (90),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (3),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                     //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                      //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                                   //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                             //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                               //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                     //          .ready
		.av_response             (),                                                                                          // (terminated)
		.av_writeresponserequest (1'b0),                                                                                      // (terminated)
		.av_writeresponsevalid   ()                                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_BEGIN_BURST           (92),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_THREAD_ID_H           (100),
		.PKT_THREAD_ID_L           (100),
		.PKT_CACHE_H               (107),
		.PKT_CACHE_L               (104),
		.PKT_DATA_SIDEBAND_H       (91),
		.PKT_DATA_SIDEBAND_L       (91),
		.PKT_QOS_H                 (93),
		.PKT_QOS_L                 (93),
		.PKT_ADDR_SIDEBAND_H       (90),
		.PKT_ADDR_SIDEBAND_L       (90),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (6),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                       //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (nios2_qsys_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                          //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (74),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.PKT_BURST_TYPE_H          (71),
		.PKT_BURST_TYPE_L          (70),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (82),
		.PKT_THREAD_ID_L           (82),
		.PKT_CACHE_H               (89),
		.PKT_CACHE_L               (86),
		.PKT_DATA_SIDEBAND_H       (73),
		.PKT_DATA_SIDEBAND_L       (73),
		.PKT_QOS_H                 (75),
		.PKT_QOS_L                 (75),
		.PKT_ADDR_SIDEBAND_H       (72),
		.PKT_ADDR_SIDEBAND_L       (72),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.ST_DATA_W                 (92),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address              (dma_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_005_src_valid),                                                 //        rp.valid
		.rp_data                 (width_adapter_005_src_data),                                                  //          .data
		.rp_channel              (width_adapter_005_src_channel),                                               //          .channel
		.rp_startofpacket        (width_adapter_005_src_startofpacket),                                         //          .startofpacket
		.rp_endofpacket          (width_adapter_005_src_endofpacket),                                           //          .endofpacket
		.rp_ready                (width_adapter_005_src_ready),                                                 //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (85),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (74),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.PKT_BURST_TYPE_H          (71),
		.PKT_BURST_TYPE_L          (70),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (82),
		.PKT_THREAD_ID_L           (82),
		.PKT_CACHE_H               (89),
		.PKT_CACHE_L               (86),
		.PKT_DATA_SIDEBAND_H       (73),
		.PKT_DATA_SIDEBAND_L       (73),
		.PKT_QOS_H                 (75),
		.PKT_QOS_L                 (75),
		.PKT_ADDR_SIDEBAND_H       (72),
		.PKT_ADDR_SIDEBAND_L       (72),
		.PKT_RESPONSE_STATUS_H     (91),
		.PKT_RESPONSE_STATUS_L     (90),
		.ST_DATA_W                 (92),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                 //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address              (dma_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_006_src_valid),                                                  //        rp.valid
		.rp_data                 (width_adapter_006_src_data),                                                   //          .data
		.rp_channel              (width_adapter_006_src_channel),                                                //          .channel
		.rp_startofpacket        (width_adapter_006_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (width_adapter_006_src_endofpacket),                                            //          .endofpacket
		.rp_ready                (width_adapter_006_src_ready),                                                  //          .ready
		.av_response             (),                                                                             // (terminated)
		.av_writeresponserequest (1'b0),                                                                         // (terminated)
		.av_writeresponsevalid   ()                                                                              // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_BEGIN_BURST           (92),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_THREAD_ID_H           (100),
		.PKT_THREAD_ID_L           (100),
		.PKT_CACHE_H               (107),
		.PKT_CACHE_L               (104),
		.PKT_DATA_SIDEBAND_H       (91),
		.PKT_DATA_SIDEBAND_L       (91),
		.PKT_QOS_H                 (93),
		.PKT_QOS_L                 (93),
		.PKT_ADDR_SIDEBAND_H       (90),
		.PKT_ADDR_SIDEBAND_L       (90),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                             //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.av_address              (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_007_src_valid),                                                              //        rp.valid
		.rp_data                 (width_adapter_007_src_data),                                                               //          .data
		.rp_channel              (width_adapter_007_src_channel),                                                            //          .channel
		.rp_startofpacket        (width_adapter_007_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (width_adapter_007_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (width_adapter_007_src_ready),                                                              //          .ready
		.av_response             (),                                                                                         // (terminated)
		.av_writeresponserequest (1'b0),                                                                                     // (terminated)
		.av_writeresponsevalid   ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (110),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (111),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (110),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                       //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                       //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                        //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                 //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                     //                .channel
		.rf_sink_ready           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (111),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (110),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                                 //                .channel
		.rf_sink_ready           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (111),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (110),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) wrapper_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (wrapper_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                 //                .channel
		.rf_sink_ready           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (111),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (255),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (344),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (287),
		.PKT_BYTEEN_L              (256),
		.PKT_ADDR_H                (319),
		.PKT_ADDR_L                (288),
		.PKT_TRANS_COMPRESSED_READ (320),
		.PKT_TRANS_POSTED          (321),
		.PKT_TRANS_WRITE           (322),
		.PKT_TRANS_READ            (323),
		.PKT_TRANS_LOCK            (324),
		.PKT_SRC_ID_H              (348),
		.PKT_SRC_ID_L              (346),
		.PKT_DEST_ID_H             (351),
		.PKT_DEST_ID_L             (349),
		.PKT_BURSTWRAP_H           (336),
		.PKT_BURSTWRAP_L           (334),
		.PKT_BYTE_CNT_H            (333),
		.PKT_BYTE_CNT_L            (326),
		.PKT_PROTECTION_H          (355),
		.PKT_PROTECTION_L          (353),
		.PKT_RESPONSE_STATUS_H     (361),
		.PKT_RESPONSE_STATUS_L     (360),
		.PKT_BURST_SIZE_H          (339),
		.PKT_BURST_SIZE_L          (337),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (362),
		.AVS_BURSTCOUNT_W          (8),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                              //                .channel
		.rf_sink_ready           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (363),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (258),
		.FIFO_DEPTH          (128),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_startofpacket  (1'b0),                                                                                // (terminated)
		.in_endofpacket    (1'b0),                                                                                // (terminated)
		.out_startofpacket (),                                                                                    // (terminated)
		.out_endofpacket   (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (110),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                  //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                  //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                   //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                            //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (111),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr2_emif_afi_clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (103),
		.PKT_PROTECTION_L          (101),
		.PKT_RESPONSE_STATUS_H     (109),
		.PKT_RESPONSE_STATUS_L     (108),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (110),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (111),
		.FIFO_DEPTH          (9),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (16),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                                          // (terminated)
		.out_startofpacket (),                                                                                              // (terminated)
		.out_endofpacket   (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_THREAD_ID_H           (71),
		.PKT_THREAD_ID_L           (71),
		.PKT_CACHE_H               (78),
		.PKT_CACHE_L               (75),
		.PKT_DATA_SIDEBAND_H       (62),
		.PKT_DATA_SIDEBAND_L       (62),
		.PKT_QOS_H                 (64),
		.PKT_QOS_L                 (64),
		.PKT_ADDR_SIDEBAND_H       (61),
		.PKT_ADDR_SIDEBAND_L       (61),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent (
		.clk                     (mem_if_ddr2_emif_afi_clk_clk),                                                               //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.av_address              (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_002_rsp_src_valid),                                                                  //        rp.valid
		.rp_data                 (limiter_002_rsp_src_data),                                                                   //          .data
		.rp_channel              (limiter_002_rsp_src_channel),                                                                //          .channel
		.rp_startofpacket        (limiter_002_rsp_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket          (limiter_002_rsp_src_endofpacket),                                                            //          .endofpacket
		.rp_ready                (limiter_002_rsp_src_ready),                                                                  //          .ready
		.av_response             (),                                                                                           // (terminated)
		.av_writeresponserequest (1'b0),                                                                                       // (terminated)
		.av_writeresponsevalid   ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (button_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                          //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                          //                .valid
		.cp_data                 (crosser_002_out_data),                                                           //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                    //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                        //                .channel
		.rf_sink_ready           (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.in_data           (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                    // (terminated)
		.csr_read          (1'b0),                                                                     // (terminated)
		.csr_write         (1'b0),                                                                     // (terminated)
		.csr_readdata      (),                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                     // (terminated)
		.almost_full_data  (),                                                                         // (terminated)
		.almost_empty_data (),                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                     // (terminated)
		.out_startofpacket (),                                                                         // (terminated)
		.out_endofpacket   (),                                                                         // (terminated)
		.in_empty          (1'b0),                                                                     // (terminated)
		.out_empty         (),                                                                         // (terminated)
		.in_error          (1'b0),                                                                     // (terminated)
		.out_error         (),                                                                         // (terminated)
		.in_channel        (1'b0),                                                                     // (terminated)
		.out_channel       ()                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_003_out_ready),                                                       //              cp.ready
		.cp_valid                (crosser_003_out_valid),                                                       //                .valid
		.cp_data                 (crosser_003_out_data),                                                        //                .data
		.cp_startofpacket        (crosser_003_out_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (crosser_003_out_endofpacket),                                                 //                .endofpacket
		.cp_channel              (crosser_003_out_channel),                                                     //                .channel
		.rf_sink_ready           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                 // (terminated)
		.csr_read          (1'b0),                                                                  // (terminated)
		.csr_write         (1'b0),                                                                  // (terminated)
		.csr_readdata      (),                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                  // (terminated)
		.almost_full_data  (),                                                                      // (terminated)
		.almost_empty_data (),                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                  // (terminated)
		.out_startofpacket (),                                                                      // (terminated)
		.out_endofpacket   (),                                                                      // (terminated)
		.in_empty          (1'b0),                                                                  // (terminated)
		.out_empty         (),                                                                      // (terminated)
		.in_error          (1'b0),                                                                  // (terminated)
		.out_error         (),                                                                      // (terminated)
		.in_channel        (1'b0),                                                                  // (terminated)
		.out_channel       ()                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_004_out_ready),                                                         //              cp.ready
		.cp_valid                (crosser_004_out_valid),                                                         //                .valid
		.cp_data                 (crosser_004_out_data),                                                          //                .data
		.cp_startofpacket        (crosser_004_out_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (crosser_004_out_endofpacket),                                                   //                .endofpacket
		.cp_channel              (crosser_004_out_channel),                                                       //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_005_out_ready),                                                                    //              cp.ready
		.cp_valid                (crosser_005_out_valid),                                                                    //                .valid
		.cp_data                 (crosser_005_out_data),                                                                     //                .data
		.cp_startofpacket        (crosser_005_out_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (crosser_005_out_endofpacket),                                                              //                .endofpacket
		.cp_channel              (crosser_005_out_channel),                                                                  //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_006_out_ready),                                                                //              cp.ready
		.cp_valid                (crosser_006_out_valid),                                                                //                .valid
		.cp_data                 (crosser_006_out_data),                                                                 //                .data
		.cp_startofpacket        (crosser_006_out_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (crosser_006_out_endofpacket),                                                          //                .endofpacket
		.cp_channel              (crosser_006_out_channel),                                                              //                .channel
		.rf_sink_ready           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_startofpacket  (1'b0),                                                                           // (terminated)
		.in_endofpacket    (1'b0),                                                                           // (terminated)
		.out_startofpacket (),                                                                               // (terminated)
		.out_endofpacket   (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (74),
		.PKT_PROTECTION_L          (72),
		.PKT_RESPONSE_STATUS_H     (80),
		.PKT_RESPONSE_STATUS_L     (79),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (81),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_007_out_ready),                                                                //              cp.ready
		.cp_valid                (crosser_007_out_valid),                                                                //                .valid
		.cp_data                 (crosser_007_out_data),                                                                 //                .data
		.cp_startofpacket        (crosser_007_out_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (crosser_007_out_endofpacket),                                                          //                .endofpacket
		.cp_channel              (crosser_007_out_channel),                                                              //                .channel
		.rf_sink_ready           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (82),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_startofpacket  (1'b0),                                                                           // (terminated)
		.in_endofpacket    (1'b0),                                                                           // (terminated)
		.out_startofpacket (),                                                                               // (terminated)
		.out_endofpacket   (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	DE4_QSYS_addr_router addr_router (
		.sink_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                     //       src.ready
		.src_valid          (addr_router_src_valid),                                                                     //          .valid
		.src_data           (addr_router_src_data),                                                                      //          .data
		.src_channel        (addr_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                //          .endofpacket
	);

	DE4_QSYS_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	DE4_QSYS_addr_router_002 addr_router_002 (
		.sink_ready         (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                   //          .valid
		.src_data           (addr_router_002_src_data),                                                    //          .data
		.src_channel        (addr_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                              //          .endofpacket
	);

	DE4_QSYS_addr_router_002 addr_router_003 (
		.sink_ready         (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                    //          .valid
		.src_data           (addr_router_003_src_data),                                                     //          .data
		.src_channel        (addr_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                               //          .endofpacket
	);

	DE4_QSYS_addr_router_004 addr_router_004 (
		.sink_ready         (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ppl_mem_reader_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                                //          .valid
		.src_data           (addr_router_004_src_data),                                                                 //          .data
		.src_channel        (addr_router_004_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                           //          .endofpacket
	);

	DE4_QSYS_id_router id_router (
		.sink_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_src_valid),                                                                     //          .valid
		.src_data           (id_router_src_data),                                                                      //          .data
		.src_channel        (id_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                //          .endofpacket
	);

	DE4_QSYS_id_router id_router_001 (
		.sink_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	DE4_QSYS_id_router_002 id_router_002 (
		.sink_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                                           //          .valid
		.src_data           (id_router_002_src_data),                                                            //          .data
		.src_channel        (id_router_002_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                      //          .endofpacket
	);

	DE4_QSYS_id_router id_router_003 (
		.sink_ready         (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (wrapper_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                 //       src.ready
		.src_valid          (id_router_003_src_valid),                                                 //          .valid
		.src_data           (id_router_003_src_data),                                                  //          .data
		.src_channel        (id_router_003_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                            //          .endofpacket
	);

	DE4_QSYS_id_router_004 id_router_004 (
		.sink_ready         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mem_if_ddr2_emif_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                         //       src.ready
		.src_valid          (id_router_004_src_valid),                                                         //          .valid
		.src_data           (id_router_004_src_data),                                                          //          .data
		.src_channel        (id_router_004_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                    //          .endofpacket
	);

	DE4_QSYS_id_router_005 id_router_005 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	DE4_QSYS_id_router_005 id_router_006 (
		.sink_ready         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_clock_crossing_bridge_io_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                   //          .valid
		.src_data           (id_router_006_src_data),                                                                    //          .data
		.src_channel        (id_router_006_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                              //          .endofpacket
	);

	DE4_QSYS_addr_router_005 addr_router_005 (
		.sink_ready         (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_clock_crossing_bridge_io_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr2_emif_afi_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                                  //          .valid
		.src_data           (addr_router_005_src_data),                                                                   //          .data
		.src_channel        (addr_router_005_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                             //          .endofpacket
	);

	DE4_QSYS_id_router_007 id_router_007 (
		.sink_ready         (button_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                              //       src.ready
		.src_valid          (id_router_007_src_valid),                                              //          .valid
		.src_data           (id_router_007_src_data),                                               //          .data
		.src_channel        (id_router_007_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                         //          .endofpacket
	);

	DE4_QSYS_id_router_007 id_router_008 (
		.sink_ready         (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                           //       src.ready
		.src_valid          (id_router_008_src_valid),                                           //          .valid
		.src_data           (id_router_008_src_data),                                            //          .data
		.src_channel        (id_router_008_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                      //          .endofpacket
	);

	DE4_QSYS_id_router_007 id_router_009 (
		.sink_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                             //       src.ready
		.src_valid          (id_router_009_src_valid),                                             //          .valid
		.src_data           (id_router_009_src_data),                                              //          .data
		.src_channel        (id_router_009_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                        //          .endofpacket
	);

	DE4_QSYS_id_router_007 id_router_010 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                        //       src.ready
		.src_valid          (id_router_010_src_valid),                                                        //          .valid
		.src_data           (id_router_010_src_data),                                                         //          .data
		.src_channel        (id_router_010_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                   //          .endofpacket
	);

	DE4_QSYS_id_router_007 id_router_011 (
		.sink_ready         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                    //       src.ready
		.src_valid          (id_router_011_src_valid),                                                    //          .valid
		.src_data           (id_router_011_src_data),                                                     //          .data
		.src_channel        (id_router_011_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                               //          .endofpacket
	);

	DE4_QSYS_id_router_007 id_router_012 (
		.sink_ready         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                    //       src.ready
		.src_valid          (id_router_012_src_valid),                                                    //          .valid
		.src_data           (id_router_012_src_data),                                                     //          .data
		.src_channel        (id_router_012_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                               //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (3),
		.PIPELINED                 (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.VALID_WIDTH               (7),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (mem_if_ddr2_emif_afi_clk_clk),   //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (99),
		.PKT_DEST_ID_L             (97),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (32),
		.PIPELINED                 (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.VALID_WIDTH               (7),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (mem_if_ddr2_emif_afi_clk_clk),       //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (70),
		.PKT_DEST_ID_L             (68),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (81),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (mem_if_ddr2_emif_afi_clk_clk),       //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_005_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_005_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_005_src_data),           //          .data
		.cmd_sink_channel       (addr_router_005_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_005_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_005_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_005_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_005_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_005_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_005_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_005_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_005_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (mem_if_ddr2_emif_afi_clk_clk),        //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_src_ready),              //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (mem_if_ddr2_emif_afi_clk_clk),            //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_001_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_001_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_001_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_001_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_001_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_001_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_002 (
		.clk                   (mem_if_ddr2_emif_afi_clk_clk),            //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_003_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_003_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_003_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_003_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_003_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_003_src_ready),              //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (mem_if_ddr2_emif_afi_clk_clk),            //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_demux_001_src4_valid),           //     sink0.valid
		.sink0_data            (cmd_xbar_demux_001_src4_data),            //          .data
		.sink0_channel         (cmd_xbar_demux_001_src4_channel),         //          .channel
		.sink0_startofpacket   (cmd_xbar_demux_001_src4_startofpacket),   //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_demux_001_src4_endofpacket),     //          .endofpacket
		.sink0_ready           (cmd_xbar_demux_001_src4_ready),           //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (110),
		.ST_CHANNEL_W              (7),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_004 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (crosser_out_valid),                       //     sink0.valid
		.sink0_data            (crosser_out_data),                        //          .data
		.sink0_channel         (crosser_out_channel),                     //          .channel
		.sink0_startofpacket   (crosser_out_startofpacket),               //          .startofpacket
		.sink0_endofpacket     (crosser_out_endofpacket),                 //          .endofpacket
		.sink0_ready           (crosser_out_ready),                       //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (mem_if_ddr2_emif_afi_clk_clk),       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~mem_if_ddr2_emif_afi_reset_reset),  // reset_in0.reset
		.clk        (mem_if_ddr2_emif_afi_clk_clk),       //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	DE4_QSYS_cmd_xbar_demux cmd_xbar_demux (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),      //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //           .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //           .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_mux_004 cmd_xbar_mux_004 (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),        //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),             //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),             //          .valid
		.sink0_channel       (width_adapter_src_channel),           //          .channel
		.sink0_data          (width_adapter_src_data),              //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),       //          .endofpacket
		.sink1_ready         (width_adapter_001_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_001_src_valid),         //          .valid
		.sink1_channel       (width_adapter_001_src_channel),       //          .channel
		.sink1_data          (width_adapter_001_src_data),          //          .data
		.sink1_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_001_src_endofpacket),   //          .endofpacket
		.sink2_ready         (width_adapter_002_src_ready),         //     sink2.ready
		.sink2_valid         (width_adapter_002_src_valid),         //          .valid
		.sink2_channel       (width_adapter_002_src_channel),       //          .channel
		.sink2_data          (width_adapter_002_src_data),          //          .data
		.sink2_startofpacket (width_adapter_002_src_startofpacket), //          .startofpacket
		.sink2_endofpacket   (width_adapter_002_src_endofpacket),   //          .endofpacket
		.sink3_ready         (width_adapter_003_src_ready),         //     sink3.ready
		.sink3_valid         (width_adapter_003_src_valid),         //          .valid
		.sink3_channel       (width_adapter_003_src_channel),       //          .channel
		.sink3_data          (width_adapter_003_src_data),          //          .data
		.sink3_startofpacket (width_adapter_003_src_startofpacket), //          .startofpacket
		.sink3_endofpacket   (width_adapter_003_src_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux rsp_xbar_demux (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),      //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_004 rsp_xbar_demux_002 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_004_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_004_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_004_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_004_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_004_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_004_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_004_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_004_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_004_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_004_src3_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_003_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (width_adapter_004_src_ready),           //     sink3.ready
		.sink3_valid         (width_adapter_004_src_valid),           //          .valid
		.sink3_channel       (width_adapter_004_src_channel),         //          .channel
		.sink3_data          (width_adapter_004_src_data),            //          .data
		.sink3_startofpacket (width_adapter_004_src_startofpacket),   //          .startofpacket
		.sink3_endofpacket   (width_adapter_004_src_endofpacket),     //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_005_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (crosser_001_out_ready),                 //     sink5.ready
		.sink5_valid         (crosser_001_out_valid),                 //          .valid
		.sink5_channel       (crosser_001_out_channel),               //          .channel
		.sink5_data          (crosser_001_out_data),                  //          .data
		.sink5_startofpacket (crosser_001_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket   (crosser_001_out_endofpacket)            //          .endofpacket
	);

	DE4_QSYS_cmd_xbar_demux_005 cmd_xbar_demux_005 (
		.clk                (mem_if_ddr2_emif_afi_clk_clk),          //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_005_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_005_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_005_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_005_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_005_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_005_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_005_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_005_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_005_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_005_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_005_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_005_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_005_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_005_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_005_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_005_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_005_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_005_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_005_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_005_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_005_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_005_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_005_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_005_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_005_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_005_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_005_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_005_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_005_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_005_src5_endofpacket)    //           .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_007 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_007 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_007 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_007 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_007 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_demux_007 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	DE4_QSYS_rsp_xbar_mux_005 rsp_xbar_mux_005 (
		.clk                 (mem_if_ddr2_emif_afi_clk_clk),       //       clk.clk
		.reset               (rst_controller_reset_out_reset),     // clk_reset.reset
		.src_ready           (rsp_xbar_mux_005_src_ready),         //       src.ready
		.src_valid           (rsp_xbar_mux_005_src_valid),         //          .valid
		.src_data            (rsp_xbar_mux_005_src_data),          //          .data
		.src_channel         (rsp_xbar_mux_005_src_channel),       //          .channel
		.src_startofpacket   (rsp_xbar_mux_005_src_startofpacket), //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_005_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_008_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_008_out_valid),              //          .valid
		.sink0_channel       (crosser_008_out_channel),            //          .channel
		.sink0_data          (crosser_008_out_data),               //          .data
		.sink0_startofpacket (crosser_008_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_008_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_009_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_009_out_valid),              //          .valid
		.sink1_channel       (crosser_009_out_channel),            //          .channel
		.sink1_data          (crosser_009_out_data),               //          .data
		.sink1_startofpacket (crosser_009_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_009_out_endofpacket),        //          .endofpacket
		.sink2_ready         (crosser_010_out_ready),              //     sink2.ready
		.sink2_valid         (crosser_010_out_valid),              //          .valid
		.sink2_channel       (crosser_010_out_channel),            //          .channel
		.sink2_data          (crosser_010_out_data),               //          .data
		.sink2_startofpacket (crosser_010_out_startofpacket),      //          .startofpacket
		.sink2_endofpacket   (crosser_010_out_endofpacket),        //          .endofpacket
		.sink3_ready         (crosser_011_out_ready),              //     sink3.ready
		.sink3_valid         (crosser_011_out_valid),              //          .valid
		.sink3_channel       (crosser_011_out_channel),            //          .channel
		.sink3_data          (crosser_011_out_data),               //          .data
		.sink3_startofpacket (crosser_011_out_startofpacket),      //          .startofpacket
		.sink3_endofpacket   (crosser_011_out_endofpacket),        //          .endofpacket
		.sink4_ready         (crosser_012_out_ready),              //     sink4.ready
		.sink4_valid         (crosser_012_out_valid),              //          .valid
		.sink4_channel       (crosser_012_out_channel),            //          .channel
		.sink4_data          (crosser_012_out_data),               //          .data
		.sink4_startofpacket (crosser_012_out_startofpacket),      //          .startofpacket
		.sink4_endofpacket   (crosser_012_out_endofpacket),        //          .endofpacket
		.sink5_ready         (crosser_013_out_ready),              //     sink5.ready
		.sink5_valid         (crosser_013_out_valid),              //          .valid
		.sink5_channel       (crosser_013_out_channel),            //          .channel
		.sink5_data          (crosser_013_out_data),               //          .data
		.sink5_startofpacket (crosser_013_out_startofpacket),      //          .startofpacket
		.sink5_endofpacket   (crosser_013_out_endofpacket)         //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (84),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (87),
		.IN_PKT_BURST_SIZE_L           (85),
		.IN_PKT_RESPONSE_STATUS_H      (109),
		.IN_PKT_RESPONSE_STATUS_L      (108),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (89),
		.IN_PKT_BURST_TYPE_L           (88),
		.IN_ST_DATA_W                  (110),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (333),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (339),
		.OUT_PKT_BURST_SIZE_L          (337),
		.OUT_PKT_RESPONSE_STATUS_H     (361),
		.OUT_PKT_RESPONSE_STATUS_L     (360),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (341),
		.OUT_PKT_BURST_TYPE_L          (340),
		.OUT_ST_DATA_W                 (362),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src3_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src3_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src3_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src3_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data             (width_adapter_src_data),                //          .data
		.out_channel          (width_adapter_src_channel),             //          .channel
		.out_valid            (width_adapter_src_valid),               //          .valid
		.out_ready            (width_adapter_src_ready),               //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),       //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (63),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (66),
		.IN_PKT_BURSTWRAP_L            (64),
		.IN_PKT_BURST_SIZE_H           (69),
		.IN_PKT_BURST_SIZE_L           (67),
		.IN_PKT_RESPONSE_STATUS_H      (91),
		.IN_PKT_RESPONSE_STATUS_L      (90),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (71),
		.IN_PKT_BURST_TYPE_L           (70),
		.IN_ST_DATA_W                  (92),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (333),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (339),
		.OUT_PKT_BURST_SIZE_L          (337),
		.OUT_PKT_RESPONSE_STATUS_H     (361),
		.OUT_PKT_RESPONSE_STATUS_L     (360),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (341),
		.OUT_PKT_BURST_TYPE_L          (340),
		.OUT_ST_DATA_W                 (362),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (63),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (66),
		.IN_PKT_BURSTWRAP_L            (64),
		.IN_PKT_BURST_SIZE_H           (69),
		.IN_PKT_BURST_SIZE_L           (67),
		.IN_PKT_RESPONSE_STATUS_H      (91),
		.IN_PKT_RESPONSE_STATUS_L      (90),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (71),
		.IN_PKT_BURST_TYPE_L           (70),
		.IN_ST_DATA_W                  (92),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (333),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (339),
		.OUT_PKT_BURST_SIZE_L          (337),
		.OUT_PKT_RESPONSE_STATUS_H     (361),
		.OUT_PKT_RESPONSE_STATUS_L     (360),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (341),
		.OUT_PKT_BURST_TYPE_L          (340),
		.OUT_ST_DATA_W                 (362),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_003_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_003_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_003_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_003_src0_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (84),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (87),
		.IN_PKT_BURST_SIZE_L           (85),
		.IN_PKT_RESPONSE_STATUS_H      (109),
		.IN_PKT_RESPONSE_STATUS_L      (108),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (89),
		.IN_PKT_BURST_TYPE_L           (88),
		.IN_ST_DATA_W                  (110),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (333),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (339),
		.OUT_PKT_BURST_SIZE_L          (337),
		.OUT_PKT_RESPONSE_STATUS_H     (361),
		.OUT_PKT_RESPONSE_STATUS_L     (360),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (341),
		.OUT_PKT_BURST_TYPE_L          (340),
		.OUT_ST_DATA_W                 (362),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_003 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_004_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_004_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_004_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_004_src0_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_003_src_data),            //          .data
		.out_channel          (width_adapter_003_src_channel),         //          .channel
		.out_valid            (width_adapter_003_src_valid),           //          .valid
		.out_ready            (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (333),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (336),
		.IN_PKT_BURSTWRAP_L            (334),
		.IN_PKT_BURST_SIZE_H           (339),
		.IN_PKT_BURST_SIZE_L           (337),
		.IN_PKT_RESPONSE_STATUS_H      (361),
		.IN_PKT_RESPONSE_STATUS_L      (360),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (341),
		.IN_PKT_BURST_TYPE_L           (340),
		.IN_ST_DATA_W                  (362),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (81),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (87),
		.OUT_PKT_BURST_SIZE_L          (85),
		.OUT_PKT_RESPONSE_STATUS_H     (109),
		.OUT_PKT_RESPONSE_STATUS_L     (108),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (89),
		.OUT_PKT_BURST_TYPE_L          (88),
		.OUT_ST_DATA_W                 (110),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_004 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_004_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_004_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_004_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_004_src0_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (333),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (336),
		.IN_PKT_BURSTWRAP_L            (334),
		.IN_PKT_BURST_SIZE_H           (339),
		.IN_PKT_BURST_SIZE_L           (337),
		.IN_PKT_RESPONSE_STATUS_H      (361),
		.IN_PKT_RESPONSE_STATUS_L      (360),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (341),
		.IN_PKT_BURST_TYPE_L           (340),
		.IN_ST_DATA_W                  (362),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (63),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (69),
		.OUT_PKT_BURST_SIZE_L          (67),
		.OUT_PKT_RESPONSE_STATUS_H     (91),
		.OUT_PKT_RESPONSE_STATUS_L     (90),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (71),
		.OUT_PKT_BURST_TYPE_L          (70),
		.OUT_ST_DATA_W                 (92),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_005 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_004_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_004_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_004_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_004_src1_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (333),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (336),
		.IN_PKT_BURSTWRAP_L            (334),
		.IN_PKT_BURST_SIZE_H           (339),
		.IN_PKT_BURST_SIZE_L           (337),
		.IN_PKT_RESPONSE_STATUS_H      (361),
		.IN_PKT_RESPONSE_STATUS_L      (360),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (341),
		.IN_PKT_BURST_TYPE_L           (340),
		.IN_ST_DATA_W                  (362),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (63),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (69),
		.OUT_PKT_BURST_SIZE_L          (67),
		.OUT_PKT_RESPONSE_STATUS_H     (91),
		.OUT_PKT_RESPONSE_STATUS_L     (90),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (71),
		.OUT_PKT_BURST_TYPE_L          (70),
		.OUT_ST_DATA_W                 (92),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_006 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_004_src2_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_004_src2_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_004_src2_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_004_src2_ready),         //          .ready
		.in_data              (rsp_xbar_demux_004_src2_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (333),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (336),
		.IN_PKT_BURSTWRAP_L            (334),
		.IN_PKT_BURST_SIZE_H           (339),
		.IN_PKT_BURST_SIZE_L           (337),
		.IN_PKT_RESPONSE_STATUS_H      (361),
		.IN_PKT_RESPONSE_STATUS_L      (360),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (341),
		.IN_PKT_BURST_TYPE_L           (340),
		.IN_ST_DATA_W                  (362),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (81),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (87),
		.OUT_PKT_BURST_SIZE_L          (85),
		.OUT_PKT_RESPONSE_STATUS_H     (109),
		.OUT_PKT_RESPONSE_STATUS_L     (108),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (89),
		.OUT_PKT_BURST_TYPE_L          (88),
		.OUT_ST_DATA_W                 (110),
		.ST_CHANNEL_W                  (7),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (mem_if_ddr2_emif_afi_clk_clk),          //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_004_src3_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_004_src3_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_004_src3_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_004_src3_ready),         //          .ready
		.in_data              (rsp_xbar_demux_004_src3_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (110),
		.BITS_PER_SYMBOL     (110),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (7),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src5_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (110),
		.BITS_PER_SYMBOL     (110),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (7),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src1_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src1_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src1_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src1_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src1_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src2_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src2_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src2_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src2_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src2_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src2_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src3_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src3_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src3_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src3_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src3_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src3_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src4_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src4_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src4_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src4_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src4_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src4_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (mem_if_ddr2_emif_afi_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src5_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_008 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_007_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_007_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_007_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_007_src0_data),          //              .data
		.out_ready         (crosser_008_out_ready),                 //           out.ready
		.out_valid         (crosser_008_out_valid),                 //              .valid
		.out_startofpacket (crosser_008_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_008_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_008_out_channel),               //              .channel
		.out_data          (crosser_008_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_009 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_009_out_ready),                 //           out.ready
		.out_valid         (crosser_009_out_valid),                 //              .valid
		.out_startofpacket (crosser_009_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_009_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_009_out_channel),               //              .channel
		.out_data          (crosser_009_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_010 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_009_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_009_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_009_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_009_src0_data),          //              .data
		.out_ready         (crosser_010_out_ready),                 //           out.ready
		.out_valid         (crosser_010_out_valid),                 //              .valid
		.out_startofpacket (crosser_010_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_010_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_010_out_channel),               //              .channel
		.out_data          (crosser_010_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_011 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_010_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_010_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_010_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_010_src0_data),          //              .data
		.out_ready         (crosser_011_out_ready),                 //           out.ready
		.out_valid         (crosser_011_out_valid),                 //              .valid
		.out_startofpacket (crosser_011_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_011_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_011_out_channel),               //              .channel
		.out_data          (crosser_011_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_012 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_011_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_011_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_011_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_011_src0_data),          //              .data
		.out_ready         (crosser_012_out_ready),                 //           out.ready
		.out_valid         (crosser_012_out_valid),                 //              .valid
		.out_startofpacket (crosser_012_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_012_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_012_out_channel),               //              .channel
		.out_data          (crosser_012_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (81),
		.BITS_PER_SYMBOL     (81),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_013 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (mem_if_ddr2_emif_afi_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_013_out_ready),                 //           out.ready
		.out_valid         (crosser_013_out_valid),                 //              .valid
		.out_startofpacket (crosser_013_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_013_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_013_out_channel),               //              .channel
		.out_data          (crosser_013_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	DE4_QSYS_irq_mapper irq_mapper (
		.clk           (mem_if_ddr2_emif_afi_clk_clk),   //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (mem_if_ddr2_emif_afi_clk_clk),       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

endmodule
