library verilog;
use verilog.vl_types.all;
entity altera_conduit_bfm_0006 is
    port(
        sig_export      : inout  vl_logic
    );
end altera_conduit_bfm_0006;
