library verilog;
use verilog.vl_types.all;
entity alt_mem_ddrx_ecc_encoder_decoder_wrapper is
    generic(
        CFG_LOCAL_DATA_WIDTH: integer := 80;
        CFG_LOCAL_ADDR_WIDTH: integer := 32;
        CFG_DWIDTH_RATIO: integer := 2;
        CFG_MEM_IF_DQ_WIDTH: integer := 40;
        CFG_MEM_IF_DQS_WIDTH: integer := 5;
        CFG_ECC_CODE_WIDTH: integer := 8;
        CFG_ECC_MULTIPLES: integer := 1;
        CFG_ECC_ENC_REG : integer := 0;
        CFG_ECC_DEC_REG : integer := 0;
        CFG_ECC_DECODER_REG: integer := 0;
        CFG_ECC_RDATA_REG: integer := 0;
        CFG_PORT_WIDTH_INTERFACE_WIDTH: integer := 8;
        CFG_PORT_WIDTH_ENABLE_ECC: integer := 1;
        CFG_PORT_WIDTH_GEN_SBE: integer := 1;
        CFG_PORT_WIDTH_GEN_DBE: integer := 1;
        CFG_PORT_WIDTH_ENABLE_INTR: integer := 1;
        CFG_PORT_WIDTH_MASK_SBE_INTR: integer := 1;
        CFG_PORT_WIDTH_MASK_DBE_INTR: integer := 1;
        CFG_PORT_WIDTH_MASK_CORR_DROPPED_INTR: integer := 1;
        CFG_PORT_WIDTH_CLR_INTR: integer := 1;
        STS_PORT_WIDTH_SBE_ERROR: integer := 1;
        STS_PORT_WIDTH_DBE_ERROR: integer := 1;
        STS_PORT_WIDTH_SBE_COUNT: integer := 8;
        STS_PORT_WIDTH_DBE_COUNT: integer := 8;
        STS_PORT_WIDTH_CORR_DROP_ERROR: integer := 1;
        STS_PORT_WIDTH_CORR_DROP_COUNT: integer := 8
    );
    port(
        ctl_clk         : in     vl_logic;
        ctl_reset_n     : in     vl_logic;
        cfg_interface_width: in     vl_logic_vector;
        cfg_enable_ecc  : in     vl_logic_vector;
        cfg_gen_sbe     : in     vl_logic_vector;
        cfg_gen_dbe     : in     vl_logic_vector;
        cfg_enable_intr : in     vl_logic_vector;
        cfg_mask_sbe_intr: in     vl_logic_vector;
        cfg_mask_dbe_intr: in     vl_logic_vector;
        cfg_mask_corr_dropped_intr: in     vl_logic_vector;
        cfg_clr_intr    : in     vl_logic_vector;
        wdatap_dm       : in     vl_logic_vector;
        wdatap_data     : in     vl_logic_vector;
        wdatap_rmw_partial_data: in     vl_logic_vector;
        wdatap_rmw_correct_data: in     vl_logic_vector;
        wdatap_rmw_partial: in     vl_logic;
        wdatap_rmw_correct: in     vl_logic;
        wdatap_ecc_code : in     vl_logic_vector;
        wdatap_ecc_code_overwrite: in     vl_logic_vector;
        rdatap_rcvd_addr: in     vl_logic_vector;
        rdatap_rcvd_cmd : in     vl_logic;
        rdatap_rcvd_corr_dropped: in     vl_logic;
        afi_rdata       : in     vl_logic_vector;
        afi_rdata_valid : in     vl_logic_vector;
        ecc_rdata       : out    vl_logic_vector;
        ecc_rdata_valid : out    vl_logic;
        ecc_dm          : out    vl_logic_vector;
        ecc_wdata       : out    vl_logic_vector;
        ecc_sbe         : out    vl_logic_vector;
        ecc_dbe         : out    vl_logic_vector;
        ecc_code        : out    vl_logic_vector;
        ecc_interrupt   : out    vl_logic;
        sts_sbe_error   : out    vl_logic_vector;
        sts_dbe_error   : out    vl_logic_vector;
        sts_sbe_count   : out    vl_logic_vector;
        sts_dbe_count   : out    vl_logic_vector;
        sts_err_addr    : out    vl_logic_vector;
        sts_corr_dropped: out    vl_logic_vector;
        sts_corr_dropped_count: out    vl_logic_vector;
        sts_corr_dropped_addr: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CFG_LOCAL_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_LOCAL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_DWIDTH_RATIO : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_CODE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_MULTIPLES : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_ENC_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_DEC_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_DECODER_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECC_RDATA_REG : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_INTERFACE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_ECC : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_GEN_SBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_GEN_DBE : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_ENABLE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MASK_SBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MASK_DBE_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_MASK_CORR_DROPPED_INTR : constant is 1;
    attribute mti_svvh_generic_type of CFG_PORT_WIDTH_CLR_INTR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_SBE_ERROR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_DBE_ERROR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_SBE_COUNT : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_DBE_COUNT : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_CORR_DROP_ERROR : constant is 1;
    attribute mti_svvh_generic_type of STS_PORT_WIDTH_CORR_DROP_COUNT : constant is 1;
end alt_mem_ddrx_ecc_encoder_decoder_wrapper;
