library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_p0 is
    generic(
        DEVICE_FAMILY   : string  := "Stratix IV";
        ALTERA_ALT_MEM_IF_PHY_FAST_SIM_MODEL: integer := 1;
        OCT_TERM_CONTROL_WIDTH: integer := 14;
        MEM_IF_ADDR_WIDTH: integer := 14;
        MEM_IF_BANKADDR_WIDTH: integer := 3;
        MEM_IF_CK_WIDTH : integer := 2;
        MEM_IF_CLK_EN_WIDTH: integer := 1;
        MEM_IF_CS_WIDTH : integer := 1;
        MEM_IF_DM_WIDTH : integer := 8;
        MEM_IF_CONTROL_WIDTH: integer := 1;
        MEM_IF_DQ_WIDTH : integer := 64;
        MEM_IF_DQS_WIDTH: integer := 8;
        MEM_IF_READ_DQS_WIDTH: integer := 8;
        MEM_IF_WRITE_DQS_WIDTH: integer := 8;
        MEM_IF_ODT_WIDTH: integer := 1;
        AFI_ADDR_WIDTH  : integer := 28;
        AFI_DM_WIDTH    : integer := 32;
        AFI_BANKADDR_WIDTH: integer := 6;
        AFI_CS_WIDTH    : integer := 2;
        AFI_CLK_EN_WIDTH: integer := 2;
        AFI_CONTROL_WIDTH: integer := 2;
        AFI_ODT_WIDTH   : integer := 2;
        AFI_DQ_WIDTH    : integer := 256;
        AFI_WRITE_DQS_WIDTH: integer := 16;
        AFI_RATE_RATIO  : integer := 2;
        AFI_WLAT_WIDTH  : integer := 6;
        AFI_RLAT_WIDTH  : integer := 6;
        DLL_DELAY_CTRL_WIDTH: integer := 6;
        NUM_SUBGROUP_PER_READ_DQS: integer := 1;
        QVLD_EXTRA_FLOP_STAGES: integer := 0;
        QVLD_WR_ADDRESS_OFFSET: integer := 4;
        READ_VALID_FIFO_SIZE: integer := 16;
        READ_FIFO_SIZE  : integer := 8;
        MAX_LATENCY_COUNT_WIDTH: integer := 4;
        MAX_WRITE_LATENCY_COUNT_WIDTH: integer := 4;
        NUM_WRITE_PATH_FLOP_STAGES: integer := 0;
        NUM_WRITE_FR_CYCLE_SHIFTS: integer := 0;
        REGISTER_C2P    : string  := "false";
        NUM_AC_FR_CYCLE_SHIFTS: integer := 0;
        LDC_MEM_CK_CPS_PHASE: integer := 0;
        MR1_ODS         : integer := 0;
        MR1_RTT         : integer := 3;
        MEM_T_WL        : integer := 3;
        SEQ_BURST_COUNT_WIDTH: integer := 1;
        DLL_OFFSET_CTRL_WIDTH: integer := 6;
        MEM_CLK_FREQ    : real    := 300.000000;
        DELAY_BUFFER_MODE: string  := "HIGH";
        DQS_DELAY_CHAIN_PHASE_SETTING: integer := 2;
        DQS_PHASE_SHIFT : integer := 7200;
        DELAYED_CLOCK_PHASE_SETTING: integer := 2;
        AFI_DEBUG_INFO_WIDTH: integer := 32;
        CALIB_REG_WIDTH : integer := 8;
        TB_PROTOCOL     : string  := "DDR2";
        TB_MEM_CLK_FREQ : string  := "300.0";
        TB_RATE         : string  := "HALF";
        TB_MEM_DQ_WIDTH : string  := "64";
        TB_MEM_DQS_WIDTH: string  := "8";
        TB_PLL_DLL_MASTER: string  := "true";
        FAST_SIM_CALIBRATION: string  := "false";
        EXTRA_VFIFO_SHIFT: integer := 0
    );
    port(
        global_reset_n  : in     vl_logic;
        soft_reset_n    : in     vl_logic;
        csr_soft_reset_req: in     vl_logic;
        parallelterminationcontrol: in     vl_logic_vector;
        seriesterminationcontrol: in     vl_logic_vector;
        pll_mem_clk     : in     vl_logic;
        pll_write_clk   : in     vl_logic;
        pll_write_clk_pre_phy_clk: in     vl_logic;
        pll_addr_cmd_clk: in     vl_logic;
        pll_avl_clk     : in     vl_logic;
        pll_config_clk  : in     vl_logic;
        pll_locked      : in     vl_logic;
        dll_pll_locked  : out    vl_logic;
        dll_delayctrl   : in     vl_logic_vector;
        dll_clk         : out    vl_logic;
        afi_reset_n     : out    vl_logic;
        afi_reset_export_n: out    vl_logic;
        afi_clk         : in     vl_logic;
        afi_half_clk    : in     vl_logic;
        afi_addr        : in     vl_logic_vector;
        afi_ba          : in     vl_logic_vector;
        afi_cke         : in     vl_logic_vector;
        afi_cs_n        : in     vl_logic_vector;
        afi_ras_n       : in     vl_logic_vector;
        afi_we_n        : in     vl_logic_vector;
        afi_cas_n       : in     vl_logic_vector;
        afi_odt         : in     vl_logic_vector;
        afi_dqs_burst   : in     vl_logic_vector;
        afi_wdata       : in     vl_logic_vector;
        afi_wdata_valid : in     vl_logic_vector;
        afi_dm          : in     vl_logic_vector;
        afi_rdata       : out    vl_logic_vector;
        afi_rdata_en    : in     vl_logic_vector;
        afi_rdata_en_full: in     vl_logic_vector;
        afi_rdata_valid : out    vl_logic_vector;
        afi_cal_success : out    vl_logic;
        afi_cal_fail    : out    vl_logic;
        afi_wlat        : out    vl_logic_vector;
        afi_rlat        : out    vl_logic_vector;
        afi_mem_clk_disable: in     vl_logic_vector;
        mem_a           : out    vl_logic_vector;
        mem_ba          : out    vl_logic_vector;
        mem_ck          : out    vl_logic_vector;
        mem_ck_n        : out    vl_logic_vector;
        mem_cke         : out    vl_logic_vector;
        mem_cs_n        : out    vl_logic_vector;
        mem_dm          : out    vl_logic_vector;
        mem_ras_n       : out    vl_logic_vector;
        mem_cas_n       : out    vl_logic_vector;
        mem_we_n        : out    vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        mem_odt         : out    vl_logic_vector;
        addr_cmd_clk    : out    vl_logic;
        avl_clk         : out    vl_logic;
        scc_clk         : out    vl_logic;
        avl_reset_n     : out    vl_logic;
        scc_reset_n     : out    vl_logic;
        scc_data        : in     vl_logic;
        scc_dqs_ena     : in     vl_logic_vector;
        scc_dqs_io_ena  : in     vl_logic_vector;
        scc_dq_ena      : in     vl_logic_vector;
        scc_dm_ena      : in     vl_logic_vector;
        scc_upd         : in     vl_logic_vector(0 downto 0);
        capture_strobe_tracking: out    vl_logic_vector;
        phy_clk         : out    vl_logic;
        phy_reset_n     : out    vl_logic;
        phy_read_latency_counter: in     vl_logic_vector;
        phy_afi_wlat    : in     vl_logic_vector;
        phy_afi_rlat    : in     vl_logic_vector;
        phy_read_increment_vfifo_fr: in     vl_logic_vector;
        phy_read_increment_vfifo_hr: in     vl_logic_vector;
        phy_read_increment_vfifo_qr: in     vl_logic_vector;
        phy_reset_mem_stable: in     vl_logic;
        phy_cal_debug_info: in     vl_logic_vector;
        phy_read_fifo_reset: in     vl_logic_vector;
        phy_vfifo_rd_en_override: in     vl_logic_vector;
        phy_cal_success : in     vl_logic;
        phy_cal_fail    : in     vl_logic;
        phy_read_fifo_q : out    vl_logic_vector;
        calib_skip_steps: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of ALTERA_ALT_MEM_IF_PHY_FAST_SIM_MODEL : constant is 1;
    attribute mti_svvh_generic_type of OCT_TERM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATE_RATIO : constant is 1;
    attribute mti_svvh_generic_type of AFI_WLAT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RLAT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DLL_DELAY_CTRL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_SUBGROUP_PER_READ_DQS : constant is 1;
    attribute mti_svvh_generic_type of QVLD_EXTRA_FLOP_STAGES : constant is 1;
    attribute mti_svvh_generic_type of QVLD_WR_ADDRESS_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of READ_FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of MAX_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_WRITE_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_WRITE_PATH_FLOP_STAGES : constant is 1;
    attribute mti_svvh_generic_type of NUM_WRITE_FR_CYCLE_SHIFTS : constant is 1;
    attribute mti_svvh_generic_type of REGISTER_C2P : constant is 1;
    attribute mti_svvh_generic_type of NUM_AC_FR_CYCLE_SHIFTS : constant is 1;
    attribute mti_svvh_generic_type of LDC_MEM_CK_CPS_PHASE : constant is 1;
    attribute mti_svvh_generic_type of MR1_ODS : constant is 1;
    attribute mti_svvh_generic_type of MR1_RTT : constant is 1;
    attribute mti_svvh_generic_type of MEM_T_WL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_BURST_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DLL_OFFSET_CTRL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of DELAY_BUFFER_MODE : constant is 1;
    attribute mti_svvh_generic_type of DQS_DELAY_CHAIN_PHASE_SETTING : constant is 1;
    attribute mti_svvh_generic_type of DQS_PHASE_SHIFT : constant is 1;
    attribute mti_svvh_generic_type of DELAYED_CLOCK_PHASE_SETTING : constant is 1;
    attribute mti_svvh_generic_type of AFI_DEBUG_INFO_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CALIB_REG_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TB_PROTOCOL : constant is 1;
    attribute mti_svvh_generic_type of TB_MEM_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of TB_RATE : constant is 1;
    attribute mti_svvh_generic_type of TB_MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TB_MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TB_PLL_DLL_MASTER : constant is 1;
    attribute mti_svvh_generic_type of FAST_SIM_CALIBRATION : constant is 1;
    attribute mti_svvh_generic_type of EXTRA_VFIFO_SHIFT : constant is 1;
end DE4_QSYS_mem_if_ddr2_emif_p0;
