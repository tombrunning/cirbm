library verilog;
use verilog.vl_types.all;
entity altera_conduit_bfm_0005 is
    port(
        sig_export      : in     vl_logic
    );
end altera_conduit_bfm_0005;
