library verilog;
use verilog.vl_types.all;
entity alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en is
    generic(
        MEM_IF_CLK_EN_WIDTH: integer := 1;
        MEM_IF_CK_WIDTH : integer := 1;
        MEM_IF_BANKADDR_WIDTH: integer := 2;
        MEM_IF_ADDR_WIDTH: integer := 14;
        MEM_IF_ROW_ADDR_WIDTH: integer := 14;
        MEM_IF_COL_ADDR_WIDTH: integer := 10;
        MEM_IF_CS_WIDTH : integer := 1;
        MEM_IF_CONTROL_WIDTH: integer := 1;
        DEVICE_DEPTH    : integer := 1;
        DEVICE_WIDTH    : integer := 1;
        MEM_IF_CS_PER_RANK: integer := 1;
        MEM_IF_DQS_WIDTH: integer := 1;
        MEM_IF_DQ_WIDTH : integer := 8;
        MEM_IF_ODT_WIDTH: integer := 1;
        MEM_MIRROR_ADDRESSING_DEC: integer := 0;
        MEM_TRTP        : integer := 3;
        MEM_TRCD        : integer := 6;
        MEM_DQS_TO_CLK_CAPTURE_DELAY: integer := 100;
        MEM_CLK_TO_DQS_CAPTURE_DELAY: integer := 100000;
        MEM_REGDIMM_ENABLED: integer := 0;
        MEM_INIT_EN     : integer := 0;
        MEM_INIT_FILE   : string  := "";
        MEM_GUARANTEED_WRITE_INIT: integer := 0;
        DAT_DATA_WIDTH  : integer := 32;
        MEM_VERBOSE     : integer := 1
    );
    port(
        mem_a           : in     vl_logic_vector;
        mem_ba          : in     vl_logic_vector;
        mem_ck          : in     vl_logic_vector;
        mem_ck_n        : in     vl_logic_vector;
        mem_cke         : in     vl_logic_vector;
        mem_cs_n        : in     vl_logic_vector;
        mem_ras_n       : in     vl_logic_vector;
        mem_cas_n       : in     vl_logic_vector;
        mem_we_n        : in     vl_logic_vector;
        mem_dm          : in     vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        mem_odt         : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MEM_IF_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_BANKADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ROW_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_COL_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DEVICE_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of DEVICE_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_CS_PER_RANK : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_MIRROR_ADDRESSING_DEC : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRTP : constant is 1;
    attribute mti_svvh_generic_type of MEM_TRCD : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_TO_CLK_CAPTURE_DELAY : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_TO_DQS_CAPTURE_DELAY : constant is 1;
    attribute mti_svvh_generic_type of MEM_REGDIMM_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of MEM_INIT_EN : constant is 1;
    attribute mti_svvh_generic_type of MEM_INIT_FILE : constant is 1;
    attribute mti_svvh_generic_type of MEM_GUARANTEED_WRITE_INIT : constant is 1;
    attribute mti_svvh_generic_type of DAT_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_VERBOSE : constant is 1;
end alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en;
