library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_p0_new_io_pads is
    generic(
        DEVICE_FAMILY   : string  := "";
        REGISTER_C2P    : string  := "";
        LDC_MEM_CK_CPS_PHASE: string  := "";
        OCT_SERIES_TERM_CONTROL_WIDTH: string  := "";
        OCT_PARALLEL_TERM_CONTROL_WIDTH: string  := "";
        MEM_ADDRESS_WIDTH: string  := "";
        MEM_BANK_WIDTH  : string  := "";
        MEM_CHIP_SELECT_WIDTH: string  := "";
        MEM_CLK_EN_WIDTH: string  := "";
        MEM_CK_WIDTH    : string  := "";
        MEM_ODT_WIDTH   : string  := "";
        MEM_DQS_WIDTH   : string  := "";
        MEM_DM_WIDTH    : string  := "";
        MEM_CONTROL_WIDTH: string  := "";
        MEM_DQ_WIDTH    : string  := "";
        MEM_READ_DQS_WIDTH: string  := "";
        MEM_WRITE_DQS_WIDTH: string  := "";
        AFI_ADDRESS_WIDTH: string  := "";
        AFI_BANK_WIDTH  : string  := "";
        AFI_CHIP_SELECT_WIDTH: string  := "";
        AFI_CLK_EN_WIDTH: string  := "";
        AFI_ODT_WIDTH   : string  := "";
        AFI_DATA_MASK_WIDTH: string  := "";
        AFI_CONTROL_WIDTH: string  := "";
        AFI_DATA_WIDTH  : string  := "";
        AFI_DQS_WIDTH   : string  := "";
        AFI_RATE_RATIO  : string  := "";
        DLL_DELAY_CTRL_WIDTH: string  := "";
        DQS_ENABLE_CTRL_WIDTH: string  := "";
        ALTDQDQS_INPUT_FREQ: string  := "";
        ALTDQDQS_DELAY_CHAIN_BUFFER_MODE: string  := "";
        ALTDQDQS_DQS_PHASE_SETTING: string  := "";
        ALTDQDQS_DQS_PHASE_SHIFT: string  := "";
        ALTDQDQS_DELAYED_CLOCK_PHASE_SETTING: string  := "";
        FAST_SIM_MODEL  : string  := "";
        IS_HHP_HPS      : string  := ""
    );
    port(
        reset_n_addr_cmd_clk: in     vl_logic;
        reset_n_afi_clk : in     vl_logic;
        phy_reset_mem_stable: in     vl_logic;
        oct_ctl_rs_value: in     vl_logic_vector;
        oct_ctl_rt_value: in     vl_logic_vector;
        phy_ddio_addr_cmd_clk: in     vl_logic;
        phy_ddio_address: in     vl_logic_vector;
        phy_ddio_bank   : in     vl_logic_vector;
        phy_ddio_cs_n   : in     vl_logic_vector;
        phy_ddio_cke    : in     vl_logic_vector;
        phy_ddio_odt    : in     vl_logic_vector;
        phy_ddio_we_n   : in     vl_logic_vector;
        phy_ddio_ras_n  : in     vl_logic_vector;
        phy_ddio_cas_n  : in     vl_logic_vector;
        phy_mem_address : out    vl_logic_vector;
        phy_mem_bank    : out    vl_logic_vector;
        phy_mem_cs_n    : out    vl_logic_vector;
        phy_mem_cke     : out    vl_logic_vector;
        phy_mem_odt     : out    vl_logic_vector;
        phy_mem_we_n    : out    vl_logic_vector;
        phy_mem_ras_n   : out    vl_logic_vector;
        phy_mem_cas_n   : out    vl_logic_vector;
        pll_afi_clk     : in     vl_logic;
        pll_mem_clk     : in     vl_logic;
        pll_write_clk   : in     vl_logic;
        pll_dqs_ena_clk : in     vl_logic;
        phy_ddio_dq     : in     vl_logic_vector;
        phy_ddio_dqs_en : in     vl_logic_vector;
        phy_ddio_oct_ena: in     vl_logic_vector;
        dqs_enable_ctrl : in     vl_logic_vector;
        phy_ddio_wrdata_en: in     vl_logic_vector;
        phy_ddio_wrdata_mask: in     vl_logic_vector;
        phy_mem_dq      : inout  vl_logic_vector;
        phy_mem_dm      : out    vl_logic_vector;
        phy_mem_ck      : out    vl_logic_vector;
        phy_mem_ck_n    : out    vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        dll_phy_delayctrl: in     vl_logic_vector;
        ddio_phy_dq     : out    vl_logic_vector;
        read_capture_clk: out    vl_logic_vector;
        scc_clk         : in     vl_logic;
        scc_data        : in     vl_logic;
        scc_dqs_ena     : in     vl_logic_vector;
        scc_dqs_io_ena  : in     vl_logic_vector;
        scc_dq_ena      : in     vl_logic_vector;
        scc_dm_ena      : in     vl_logic_vector;
        scc_sr_dqsenable_delayctrl: in     vl_logic_vector(7 downto 0);
        scc_sr_dqsdisablen_delayctrl: in     vl_logic_vector(7 downto 0);
        scc_sr_multirank_delayctrl: in     vl_logic_vector(7 downto 0);
        scc_upd         : in     vl_logic_vector(0 downto 0);
        enable_mem_clk  : in     vl_logic_vector;
        capture_strobe_tracking: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of REGISTER_C2P : constant is 1;
    attribute mti_svvh_generic_type of LDC_MEM_CK_CPS_PHASE : constant is 1;
    attribute mti_svvh_generic_type of OCT_SERIES_TERM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of OCT_PARALLEL_TERM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CHIP_SELECT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CHIP_SELECT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DATA_MASK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATE_RATIO : constant is 1;
    attribute mti_svvh_generic_type of DLL_DELAY_CTRL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DQS_ENABLE_CTRL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_INPUT_FREQ : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DELAY_CHAIN_BUFFER_MODE : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DQS_PHASE_SETTING : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DQS_PHASE_SHIFT : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DELAYED_CLOCK_PHASE_SETTING : constant is 1;
    attribute mti_svvh_generic_type of FAST_SIM_MODEL : constant is 1;
    attribute mti_svvh_generic_type of IS_HHP_HPS : constant is 1;
end DE4_QSYS_mem_if_ddr2_emif_p0_new_io_pads;
