library verilog;
use verilog.vl_types.all;
entity DE4_QSYS_mem_if_ddr2_emif_p0_memphy is
    generic(
        DEVICE_FAMILY   : string  := "";
        OCT_SERIES_TERM_CONTROL_WIDTH: string  := "";
        OCT_PARALLEL_TERM_CONTROL_WIDTH: string  := "";
        MEM_ADDRESS_WIDTH: string  := "";
        MEM_BANK_WIDTH  : string  := "";
        MEM_CLK_EN_WIDTH: string  := "";
        MEM_CK_WIDTH    : string  := "";
        MEM_ODT_WIDTH   : string  := "";
        MEM_DQS_WIDTH   : string  := "";
        MEM_CHIP_SELECT_WIDTH: string  := "";
        MEM_CONTROL_WIDTH: string  := "";
        MEM_DM_WIDTH    : string  := "";
        MEM_DQ_WIDTH    : string  := "";
        MEM_READ_DQS_WIDTH: string  := "";
        MEM_WRITE_DQS_WIDTH: string  := "";
        MEM_IF_NUMBER_OF_RANKS: string  := "";
        AFI_ADDRESS_WIDTH: string  := "";
        AFI_DEBUG_INFO_WIDTH: string  := "";
        AFI_BANK_WIDTH  : string  := "";
        AFI_CHIP_SELECT_WIDTH: string  := "";
        AFI_CLK_EN_WIDTH: string  := "";
        AFI_ODT_WIDTH   : string  := "";
        AFI_MAX_WRITE_LATENCY_COUNT_WIDTH: string  := "";
        AFI_MAX_READ_LATENCY_COUNT_WIDTH: string  := "";
        AFI_DATA_MASK_WIDTH: string  := "";
        AFI_CONTROL_WIDTH: string  := "";
        AFI_DATA_WIDTH  : string  := "";
        AFI_DQS_WIDTH   : string  := "";
        AFI_RATE_RATIO  : string  := "";
        AFI_RRANK_WIDTH : string  := "";
        AFI_WRANK_WIDTH : string  := "";
        DLL_DELAY_CTRL_WIDTH: string  := "";
        NUM_SUBGROUP_PER_READ_DQS: string  := "";
        QVLD_EXTRA_FLOP_STAGES: string  := "";
        QVLD_WR_ADDRESS_OFFSET: string  := "";
        READ_VALID_FIFO_SIZE: string  := "";
        READ_FIFO_SIZE  : string  := "";
        MAX_LATENCY_COUNT_WIDTH: string  := "";
        MAX_READ_LATENCY: string  := "";
        MAX_WRITE_LATENCY_COUNT_WIDTH: string  := "";
        NUM_WRITE_PATH_FLOP_STAGES: string  := "";
        NUM_WRITE_FR_CYCLE_SHIFTS: string  := "";
        REGISTER_C2P    : string  := "";
        LDC_MEM_CK_CPS_PHASE: string  := "";
        NUM_AC_FR_CYCLE_SHIFTS: string  := "";
        MEM_T_RL        : string  := "";
        MR1_ODS         : string  := "";
        MR1_RTT         : string  := "";
        ALTDQDQS_INPUT_FREQ: string  := "";
        ALTDQDQS_DELAY_CHAIN_BUFFER_MODE: string  := "";
        ALTDQDQS_DQS_PHASE_SETTING: string  := "";
        ALTDQDQS_DQS_PHASE_SHIFT: string  := "";
        ALTDQDQS_DELAYED_CLOCK_PHASE_SETTING: string  := "";
        EXTRA_VFIFO_SHIFT: integer := 0;
        TB_PROTOCOL     : string  := "";
        TB_MEM_CLK_FREQ : string  := "";
        TB_RATE         : string  := "";
        TB_MEM_DQ_WIDTH : string  := "";
        TB_MEM_DQS_WIDTH: string  := "";
        TB_PLL_DLL_MASTER: string  := "";
        FAST_SIM_MODEL  : string  := "";
        FAST_SIM_CALIBRATION: string  := "";
        CALIB_REG_WIDTH : string  := ""
    );
    port(
        global_reset_n  : in     vl_logic;
        soft_reset_n    : in     vl_logic;
        ctl_reset_n     : out    vl_logic;
        ctl_reset_export_n: out    vl_logic;
        pll_locked      : in     vl_logic;
        oct_ctl_rs_value: in     vl_logic_vector;
        oct_ctl_rt_value: in     vl_logic_vector;
        afi_addr        : in     vl_logic_vector;
        afi_cke         : in     vl_logic_vector;
        afi_cs_n        : in     vl_logic_vector;
        afi_ba          : in     vl_logic_vector;
        afi_cas_n       : in     vl_logic_vector;
        afi_odt         : in     vl_logic_vector;
        afi_ras_n       : in     vl_logic_vector;
        afi_we_n        : in     vl_logic_vector;
        afi_mem_clk_disable: in     vl_logic_vector;
        afi_dqs_burst   : in     vl_logic_vector;
        afi_wlat        : out    vl_logic_vector;
        afi_rlat        : out    vl_logic_vector;
        afi_wdata       : in     vl_logic_vector;
        afi_wdata_valid : in     vl_logic_vector;
        afi_dm          : in     vl_logic_vector;
        afi_rdata       : out    vl_logic_vector;
        afi_rdata_en    : in     vl_logic_vector;
        afi_rdata_en_full: in     vl_logic_vector;
        afi_rdata_valid : out    vl_logic_vector;
        afi_cal_debug_info: out    vl_logic_vector;
        afi_cal_success : in     vl_logic;
        afi_cal_fail    : in     vl_logic;
        mem_a           : out    vl_logic_vector;
        mem_ba          : out    vl_logic_vector;
        mem_ck          : out    vl_logic_vector;
        mem_ck_n        : out    vl_logic_vector;
        mem_cke         : out    vl_logic_vector;
        mem_cs_n        : out    vl_logic_vector;
        mem_dm          : out    vl_logic_vector;
        mem_odt         : out    vl_logic_vector;
        mem_ras_n       : out    vl_logic_vector;
        mem_cas_n       : out    vl_logic_vector;
        mem_we_n        : out    vl_logic_vector;
        mem_dq          : inout  vl_logic_vector;
        mem_dqs         : inout  vl_logic_vector;
        mem_dqs_n       : inout  vl_logic_vector;
        reset_n_scc_clk : out    vl_logic;
        reset_n_avl_clk : out    vl_logic;
        scc_data        : in     vl_logic;
        scc_dqs_ena     : in     vl_logic_vector;
        scc_dqs_io_ena  : in     vl_logic_vector;
        scc_dq_ena      : in     vl_logic_vector;
        scc_dm_ena      : in     vl_logic_vector;
        scc_upd         : in     vl_logic_vector(0 downto 0);
        scc_sr_dqsenable_delayctrl: in     vl_logic_vector(7 downto 0);
        scc_sr_dqsdisablen_delayctrl: in     vl_logic_vector(7 downto 0);
        scc_sr_multirank_delayctrl: in     vl_logic_vector(7 downto 0);
        capture_strobe_tracking: out    vl_logic_vector;
        phy_clk         : out    vl_logic;
        phy_reset_n     : out    vl_logic;
        phy_read_latency_counter: in     vl_logic_vector;
        phy_afi_wlat    : in     vl_logic_vector;
        phy_afi_rlat    : in     vl_logic_vector;
        phy_num_write_fr_cycle_shifts: in     vl_logic_vector;
        phy_read_increment_vfifo_fr: in     vl_logic_vector;
        phy_read_increment_vfifo_hr: in     vl_logic_vector;
        phy_read_increment_vfifo_qr: in     vl_logic_vector;
        phy_reset_mem_stable: in     vl_logic;
        phy_cal_debug_info: in     vl_logic_vector;
        phy_read_fifo_reset: in     vl_logic_vector;
        phy_vfifo_rd_en_override: in     vl_logic_vector;
        phy_read_fifo_q : out    vl_logic_vector;
        calib_skip_steps: out    vl_logic_vector;
        pll_afi_clk     : in     vl_logic;
        pll_afi_half_clk: in     vl_logic;
        pll_addr_cmd_clk: in     vl_logic;
        pll_mem_clk     : in     vl_logic;
        pll_write_clk   : in     vl_logic;
        pll_write_clk_pre_phy_clk: in     vl_logic;
        pll_dqs_ena_clk : in     vl_logic;
        seq_clk         : in     vl_logic;
        pll_avl_clk     : in     vl_logic;
        pll_config_clk  : in     vl_logic;
        dll_clk         : out    vl_logic;
        dll_pll_locked  : out    vl_logic;
        dll_phy_delayctrl: in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DEVICE_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of OCT_SERIES_TERM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of OCT_PARALLEL_TERM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CHIP_SELECT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DM_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_READ_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_WRITE_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MEM_IF_NUMBER_OF_RANKS : constant is 1;
    attribute mti_svvh_generic_type of AFI_ADDRESS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DEBUG_INFO_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_BANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CHIP_SELECT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CLK_EN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_ODT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_MAX_WRITE_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_MAX_READ_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DATA_MASK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_CONTROL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_RATE_RATIO : constant is 1;
    attribute mti_svvh_generic_type of AFI_RRANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of AFI_WRANK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DLL_DELAY_CTRL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_SUBGROUP_PER_READ_DQS : constant is 1;
    attribute mti_svvh_generic_type of QVLD_EXTRA_FLOP_STAGES : constant is 1;
    attribute mti_svvh_generic_type of QVLD_WR_ADDRESS_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of READ_VALID_FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of READ_FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of MAX_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MAX_READ_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of MAX_WRITE_LATENCY_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_WRITE_PATH_FLOP_STAGES : constant is 1;
    attribute mti_svvh_generic_type of NUM_WRITE_FR_CYCLE_SHIFTS : constant is 1;
    attribute mti_svvh_generic_type of REGISTER_C2P : constant is 1;
    attribute mti_svvh_generic_type of LDC_MEM_CK_CPS_PHASE : constant is 1;
    attribute mti_svvh_generic_type of NUM_AC_FR_CYCLE_SHIFTS : constant is 1;
    attribute mti_svvh_generic_type of MEM_T_RL : constant is 1;
    attribute mti_svvh_generic_type of MR1_ODS : constant is 1;
    attribute mti_svvh_generic_type of MR1_RTT : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_INPUT_FREQ : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DELAY_CHAIN_BUFFER_MODE : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DQS_PHASE_SETTING : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DQS_PHASE_SHIFT : constant is 1;
    attribute mti_svvh_generic_type of ALTDQDQS_DELAYED_CLOCK_PHASE_SETTING : constant is 1;
    attribute mti_svvh_generic_type of EXTRA_VFIFO_SHIFT : constant is 1;
    attribute mti_svvh_generic_type of TB_PROTOCOL : constant is 1;
    attribute mti_svvh_generic_type of TB_MEM_CLK_FREQ : constant is 1;
    attribute mti_svvh_generic_type of TB_RATE : constant is 1;
    attribute mti_svvh_generic_type of TB_MEM_DQ_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TB_MEM_DQS_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of TB_PLL_DLL_MASTER : constant is 1;
    attribute mti_svvh_generic_type of FAST_SIM_MODEL : constant is 1;
    attribute mti_svvh_generic_type of FAST_SIM_CALIBRATION : constant is 1;
    attribute mti_svvh_generic_type of CALIB_REG_WIDTH : constant is 1;
end DE4_QSYS_mem_if_ddr2_emif_p0_memphy;
